/*
ascii码取模
注意！由于从空格开始取模，故在ascii码的基础上减去32才可正确调用
*/
`timescale 1 ns / 100 ps
module char_ram (address, q);

    input wire [11:0] address;
    output reg [7:0] q;
	 
	always @ (*)
		case(address)
			12'h000: q = 8'h00;
            12'h001: q = 8'h00;
            12'h002: q = 8'h00;
            12'h003: q = 8'h00;
            12'h004: q = 8'h00;
            12'h005: q = 8'h00;
            12'h006: q = 8'h00;
            12'h007: q = 8'h00;
            12'h008: q = 8'h00;
            12'h009: q = 8'h00;
            12'h00A: q = 8'h00;
            12'h00B: q = 8'h00;
            12'h00C: q = 8'h00;
            12'h00D: q = 8'h00;
            12'h00E: q = 8'h04;
            12'h00F: q = 8'h04;
            12'h010: q = 8'h04;
            12'h011: q = 8'h04;
            12'h012: q = 8'h04;
            12'h013: q = 8'h04;
            12'h014: q = 8'h00;
            12'h015: q = 8'h04;
            12'h016: q = 8'h00;
            12'h017: q = 8'h00;
            12'h018: q = 8'h00;
            12'h019: q = 8'h14;
            12'h01A: q = 8'h0A;
            12'h01B: q = 8'h0A;
            12'h01C: q = 8'h00;
            12'h01D: q = 8'h00;
            12'h01E: q = 8'h00;
            12'h01F: q = 8'h00;
            12'h020: q = 8'h00;
            12'h021: q = 8'h00;
            12'h022: q = 8'h00;
            12'h023: q = 8'h00;
            12'h024: q = 8'h00;
            12'h025: q = 8'h00;
            12'h026: q = 8'h14;
            12'h027: q = 8'h14;
            12'h028: q = 8'h3F;
            12'h029: q = 8'h14;
            12'h02A: q = 8'h0A;
            12'h02B: q = 8'h3F;
            12'h02C: q = 8'h0A;
            12'h02D: q = 8'h0A;
            12'h02E: q = 8'h00;
            12'h02F: q = 8'h00;
            12'h030: q = 8'h00;
            12'h031: q = 8'h04;
            12'h032: q = 8'h1E;
            12'h033: q = 8'h15;
            12'h034: q = 8'h05;
            12'h035: q = 8'h06;
            12'h036: q = 8'h0C;
            12'h037: q = 8'h14;
            12'h038: q = 8'h15;
            12'h039: q = 8'h0F;
            12'h03A: q = 8'h04;
            12'h03B: q = 8'h00;
            12'h03C: q = 8'h00;
            12'h03D: q = 8'h00;
            12'h03E: q = 8'h12;
            12'h03F: q = 8'h15;
            12'h040: q = 8'h0D;
            12'h041: q = 8'h0A;
            12'h042: q = 8'h14;
            12'h043: q = 8'h2C;
            12'h044: q = 8'h2A;
            12'h045: q = 8'h12;
            12'h046: q = 8'h00;
            12'h047: q = 8'h00;
            12'h048: q = 8'h00;
            12'h049: q = 8'h00;
            12'h04A: q = 8'h04;
            12'h04B: q = 8'h0A;
            12'h04C: q = 8'h0A;
            12'h04D: q = 8'h1E;
            12'h04E: q = 8'h15;
            12'h04F: q = 8'h15;
            12'h050: q = 8'h09;
            12'h051: q = 8'h36;
            12'h052: q = 8'h00;
            12'h053: q = 8'h00;
            12'h054: q = 8'h00;
            12'h055: q = 8'h02;
            12'h056: q = 8'h02;
            12'h057: q = 8'h01;
            12'h058: q = 8'h00;
            12'h059: q = 8'h00;
            12'h05A: q = 8'h00;
            12'h05B: q = 8'h00;
            12'h05C: q = 8'h00;
            12'h05D: q = 8'h00;
            12'h05E: q = 8'h00;
            12'h05F: q = 8'h00;
            12'h060: q = 8'h00;
            12'h061: q = 8'h20;
            12'h062: q = 8'h10;
            12'h063: q = 8'h08;
            12'h064: q = 8'h08;
            12'h065: q = 8'h08;
            12'h066: q = 8'h08;
            12'h067: q = 8'h08;
            12'h068: q = 8'h08;
            12'h069: q = 8'h10;
            12'h06A: q = 8'h20;
            12'h06B: q = 8'h00;
            12'h06C: q = 8'h00;
            12'h06D: q = 8'h02;
            12'h06E: q = 8'h04;
            12'h06F: q = 8'h08;
            12'h070: q = 8'h08;
            12'h071: q = 8'h08;
            12'h072: q = 8'h08;
            12'h073: q = 8'h08;
            12'h074: q = 8'h08;
            12'h075: q = 8'h04;
            12'h076: q = 8'h02;
            12'h077: q = 8'h00;
            12'h078: q = 8'h00;
            12'h079: q = 8'h00;
            12'h07A: q = 8'h00;
            12'h07B: q = 8'h04;
            12'h07C: q = 8'h15;
            12'h07D: q = 8'h0E;
            12'h07E: q = 8'h0E;
            12'h07F: q = 8'h15;
            12'h080: q = 8'h04;
            12'h081: q = 8'h00;
            12'h082: q = 8'h00;
            12'h083: q = 8'h00;
            12'h084: q = 8'h00;
            12'h085: q = 8'h00;
            12'h086: q = 8'h04;
            12'h087: q = 8'h04;
            12'h088: q = 8'h04;
            12'h089: q = 8'h1F;
            12'h08A: q = 8'h04;
            12'h08B: q = 8'h04;
            12'h08C: q = 8'h04;
            12'h08D: q = 8'h00;
            12'h08E: q = 8'h00;
            12'h08F: q = 8'h00;
            12'h090: q = 8'h00;
            12'h091: q = 8'h00;
            12'h092: q = 8'h00;
            12'h093: q = 8'h00;
            12'h094: q = 8'h00;
            12'h095: q = 8'h00;
            12'h096: q = 8'h00;
            12'h097: q = 8'h00;
            12'h098: q = 8'h00;
            12'h099: q = 8'h02;
            12'h09A: q = 8'h02;
            12'h09B: q = 8'h01;
            12'h09C: q = 8'h00;
            12'h09D: q = 8'h00;
            12'h09E: q = 8'h00;
            12'h09F: q = 8'h00;
            12'h0A0: q = 8'h00;
            12'h0A1: q = 8'h1F;
            12'h0A2: q = 8'h00;
            12'h0A3: q = 8'h00;
            12'h0A4: q = 8'h00;
            12'h0A5: q = 8'h00;
            12'h0A6: q = 8'h00;
            12'h0A7: q = 8'h00;
            12'h0A8: q = 8'h00;
            12'h0A9: q = 8'h00;
            12'h0AA: q = 8'h00;
            12'h0AB: q = 8'h00;
            12'h0AC: q = 8'h00;
            12'h0AD: q = 8'h00;
            12'h0AE: q = 8'h00;
            12'h0AF: q = 8'h00;
            12'h0B0: q = 8'h00;
            12'h0B1: q = 8'h02;
            12'h0B2: q = 8'h00;
            12'h0B3: q = 8'h00;
            12'h0B4: q = 8'h00;
            12'h0B5: q = 8'h10;
            12'h0B6: q = 8'h08;
            12'h0B7: q = 8'h08;
            12'h0B8: q = 8'h08;
            12'h0B9: q = 8'h04;
            12'h0BA: q = 8'h04;
            12'h0BB: q = 8'h02;
            12'h0BC: q = 8'h02;
            12'h0BD: q = 8'h02;
            12'h0BE: q = 8'h01;
            12'h0BF: q = 8'h00;
            12'h0C0: q = 8'h00;
            12'h0C1: q = 8'h00;
            12'h0C2: q = 8'h0E;
            12'h0C3: q = 8'h11;
            12'h0C4: q = 8'h11;
            12'h0C5: q = 8'h11;
            12'h0C6: q = 8'h11;
            12'h0C7: q = 8'h11;
            12'h0C8: q = 8'h11;
            12'h0C9: q = 8'h0E;
            12'h0CA: q = 8'h00;
            12'h0CB: q = 8'h00;
            12'h0CC: q = 8'h00;
            12'h0CD: q = 8'h00;
            12'h0CE: q = 8'h04;
            12'h0CF: q = 8'h06;
            12'h0D0: q = 8'h04;
            12'h0D1: q = 8'h04;
            12'h0D2: q = 8'h04;
            12'h0D3: q = 8'h04;
            12'h0D4: q = 8'h04;
            12'h0D5: q = 8'h0E;
            12'h0D6: q = 8'h00;
            12'h0D7: q = 8'h00;
            12'h0D8: q = 8'h00;
            12'h0D9: q = 8'h00;
            12'h0DA: q = 8'h0E;
            12'h0DB: q = 8'h11;
            12'h0DC: q = 8'h11;
            12'h0DD: q = 8'h08;
            12'h0DE: q = 8'h04;
            12'h0DF: q = 8'h02;
            12'h0E0: q = 8'h01;
            12'h0E1: q = 8'h1F;
            12'h0E2: q = 8'h00;
            12'h0E3: q = 8'h00;
            12'h0E4: q = 8'h00;
            12'h0E5: q = 8'h00;
            12'h0E6: q = 8'h0E;
            12'h0E7: q = 8'h11;
            12'h0E8: q = 8'h10;
            12'h0E9: q = 8'h0C;
            12'h0EA: q = 8'h10;
            12'h0EB: q = 8'h10;
            12'h0EC: q = 8'h11;
            12'h0ED: q = 8'h0E;
            12'h0EE: q = 8'h00;
            12'h0EF: q = 8'h00;
            12'h0F0: q = 8'h00;
            12'h0F1: q = 8'h00;
            12'h0F2: q = 8'h08;
            12'h0F3: q = 8'h0C;
            12'h0F4: q = 8'h0A;
            12'h0F5: q = 8'h0A;
            12'h0F6: q = 8'h09;
            12'h0F7: q = 8'h1E;
            12'h0F8: q = 8'h08;
            12'h0F9: q = 8'h18;
            12'h0FA: q = 8'h00;
            12'h0FB: q = 8'h00;
            12'h0FC: q = 8'h00;
            12'h0FD: q = 8'h00;
            12'h0FE: q = 8'h1F;
            12'h0FF: q = 8'h01;
            12'h100: q = 8'h01;
            12'h101: q = 8'h0F;
            12'h102: q = 8'h10;
            12'h103: q = 8'h10;
            12'h104: q = 8'h11;
            12'h105: q = 8'h0E;
            12'h106: q = 8'h00;
            12'h107: q = 8'h00;
            12'h108: q = 8'h00;
            12'h109: q = 8'h00;
            12'h10A: q = 8'h0E;
            12'h10B: q = 8'h09;
            12'h10C: q = 8'h01;
            12'h10D: q = 8'h0F;
            12'h10E: q = 8'h11;
            12'h10F: q = 8'h11;
            12'h110: q = 8'h11;
            12'h111: q = 8'h0E;
            12'h112: q = 8'h00;
            12'h113: q = 8'h00;
            12'h114: q = 8'h00;
            12'h115: q = 8'h00;
            12'h116: q = 8'h1F;
            12'h117: q = 8'h09;
            12'h118: q = 8'h08;
            12'h119: q = 8'h04;
            12'h11A: q = 8'h04;
            12'h11B: q = 8'h04;
            12'h11C: q = 8'h04;
            12'h11D: q = 8'h04;
            12'h11E: q = 8'h00;
            12'h11F: q = 8'h00;
            12'h120: q = 8'h00;
            12'h121: q = 8'h00;
            12'h122: q = 8'h0E;
            12'h123: q = 8'h11;
            12'h124: q = 8'h11;
            12'h125: q = 8'h0E;
            12'h126: q = 8'h11;
            12'h127: q = 8'h11;
            12'h128: q = 8'h11;
            12'h129: q = 8'h0E;
            12'h12A: q = 8'h00;
            12'h12B: q = 8'h00;
            12'h12C: q = 8'h00;
            12'h12D: q = 8'h00;
            12'h12E: q = 8'h0E;
            12'h12F: q = 8'h11;
            12'h130: q = 8'h11;
            12'h131: q = 8'h11;
            12'h132: q = 8'h1E;
            12'h133: q = 8'h10;
            12'h134: q = 8'h12;
            12'h135: q = 8'h0E;
            12'h136: q = 8'h00;
            12'h137: q = 8'h00;
            12'h138: q = 8'h00;
            12'h139: q = 8'h00;
            12'h13A: q = 8'h00;
            12'h13B: q = 8'h00;
            12'h13C: q = 8'h04;
            12'h13D: q = 8'h00;
            12'h13E: q = 8'h00;
            12'h13F: q = 8'h00;
            12'h140: q = 8'h00;
            12'h141: q = 8'h04;
            12'h142: q = 8'h00;
            12'h143: q = 8'h00;
            12'h144: q = 8'h00;
            12'h145: q = 8'h00;
            12'h146: q = 8'h00;
            12'h147: q = 8'h00;
            12'h148: q = 8'h00;
            12'h149: q = 8'h04;
            12'h14A: q = 8'h00;
            12'h14B: q = 8'h00;
            12'h14C: q = 8'h00;
            12'h14D: q = 8'h04;
            12'h14E: q = 8'h04;
            12'h14F: q = 8'h00;
            12'h150: q = 8'h00;
            12'h151: q = 8'h20;
            12'h152: q = 8'h10;
            12'h153: q = 8'h08;
            12'h154: q = 8'h04;
            12'h155: q = 8'h02;
            12'h156: q = 8'h04;
            12'h157: q = 8'h08;
            12'h158: q = 8'h10;
            12'h159: q = 8'h20;
            12'h15A: q = 8'h00;
            12'h15B: q = 8'h00;
            12'h15C: q = 8'h00;
            12'h15D: q = 8'h00;
            12'h15E: q = 8'h00;
            12'h15F: q = 8'h00;
            12'h160: q = 8'h1F;
            12'h161: q = 8'h00;
            12'h162: q = 8'h00;
            12'h163: q = 8'h1F;
            12'h164: q = 8'h00;
            12'h165: q = 8'h00;
            12'h166: q = 8'h00;
            12'h167: q = 8'h00;
            12'h168: q = 8'h00;
            12'h169: q = 8'h02;
            12'h16A: q = 8'h04;
            12'h16B: q = 8'h08;
            12'h16C: q = 8'h10;
            12'h16D: q = 8'h20;
            12'h16E: q = 8'h10;
            12'h16F: q = 8'h08;
            12'h170: q = 8'h04;
            12'h171: q = 8'h02;
            12'h172: q = 8'h00;
            12'h173: q = 8'h00;
            12'h174: q = 8'h00;
            12'h175: q = 8'h00;
            12'h176: q = 8'h0E;
            12'h177: q = 8'h11;
            12'h178: q = 8'h11;
            12'h179: q = 8'h08;
            12'h17A: q = 8'h04;
            12'h17B: q = 8'h04;
            12'h17C: q = 8'h00;
            12'h17D: q = 8'h04;
            12'h17E: q = 8'h00;
            12'h17F: q = 8'h00;
            12'h180: q = 8'h00;
            12'h181: q = 8'h00;
            12'h182: q = 8'h0E;
            12'h183: q = 8'h11;
            12'h184: q = 8'h19;
            12'h185: q = 8'h15;
            12'h186: q = 8'h15;
            12'h187: q = 8'h1D;
            12'h188: q = 8'h01;
            12'h189: q = 8'h1E;
            12'h18A: q = 8'h00;
            12'h18B: q = 8'h00;
            12'h18C: q = 8'h00;
            12'h18D: q = 8'h00;
            12'h18E: q = 8'h04;
            12'h18F: q = 8'h04;
            12'h190: q = 8'h0C;
            12'h191: q = 8'h0A;
            12'h192: q = 8'h0A;
            12'h193: q = 8'h1E;
            12'h194: q = 8'h12;
            12'h195: q = 8'h33;
            12'h196: q = 8'h00;
            12'h197: q = 8'h00;
            12'h198: q = 8'h00;
            12'h199: q = 8'h00;
            12'h19A: q = 8'h0F;
            12'h19B: q = 8'h12;
            12'h19C: q = 8'h12;
            12'h19D: q = 8'h0E;
            12'h19E: q = 8'h12;
            12'h19F: q = 8'h12;
            12'h1A0: q = 8'h12;
            12'h1A1: q = 8'h0F;
            12'h1A2: q = 8'h00;
            12'h1A3: q = 8'h00;
            12'h1A4: q = 8'h00;
            12'h1A5: q = 8'h00;
            12'h1A6: q = 8'h1E;
            12'h1A7: q = 8'h11;
            12'h1A8: q = 8'h01;
            12'h1A9: q = 8'h01;
            12'h1AA: q = 8'h01;
            12'h1AB: q = 8'h01;
            12'h1AC: q = 8'h11;
            12'h1AD: q = 8'h0E;
            12'h1AE: q = 8'h00;
            12'h1AF: q = 8'h00;
            12'h1B0: q = 8'h00;
            12'h1B1: q = 8'h00;
            12'h1B2: q = 8'h0F;
            12'h1B3: q = 8'h12;
            12'h1B4: q = 8'h12;
            12'h1B5: q = 8'h12;
            12'h1B6: q = 8'h12;
            12'h1B7: q = 8'h12;
            12'h1B8: q = 8'h12;
            12'h1B9: q = 8'h0F;
            12'h1BA: q = 8'h00;
            12'h1BB: q = 8'h00;
            12'h1BC: q = 8'h00;
            12'h1BD: q = 8'h00;
            12'h1BE: q = 8'h1F;
            12'h1BF: q = 8'h12;
            12'h1C0: q = 8'h0A;
            12'h1C1: q = 8'h0E;
            12'h1C2: q = 8'h0A;
            12'h1C3: q = 8'h02;
            12'h1C4: q = 8'h12;
            12'h1C5: q = 8'h1F;
            12'h1C6: q = 8'h00;
            12'h1C7: q = 8'h00;
            12'h1C8: q = 8'h00;
            12'h1C9: q = 8'h00;
            12'h1CA: q = 8'h1F;
            12'h1CB: q = 8'h12;
            12'h1CC: q = 8'h0A;
            12'h1CD: q = 8'h0E;
            12'h1CE: q = 8'h0A;
            12'h1CF: q = 8'h02;
            12'h1D0: q = 8'h02;
            12'h1D1: q = 8'h07;
            12'h1D2: q = 8'h00;
            12'h1D3: q = 8'h00;
            12'h1D4: q = 8'h00;
            12'h1D5: q = 8'h00;
            12'h1D6: q = 8'h1C;
            12'h1D7: q = 8'h12;
            12'h1D8: q = 8'h01;
            12'h1D9: q = 8'h01;
            12'h1DA: q = 8'h39;
            12'h1DB: q = 8'h11;
            12'h1DC: q = 8'h12;
            12'h1DD: q = 8'h0C;
            12'h1DE: q = 8'h00;
            12'h1DF: q = 8'h00;
            12'h1E0: q = 8'h00;
            12'h1E1: q = 8'h00;
            12'h1E2: q = 8'h33;
            12'h1E3: q = 8'h12;
            12'h1E4: q = 8'h12;
            12'h1E5: q = 8'h1E;
            12'h1E6: q = 8'h12;
            12'h1E7: q = 8'h12;
            12'h1E8: q = 8'h12;
            12'h1E9: q = 8'h33;
            12'h1EA: q = 8'h00;
            12'h1EB: q = 8'h00;
            12'h1EC: q = 8'h00;
            12'h1ED: q = 8'h00;
            12'h1EE: q = 8'h1F;
            12'h1EF: q = 8'h04;
            12'h1F0: q = 8'h04;
            12'h1F1: q = 8'h04;
            12'h1F2: q = 8'h04;
            12'h1F3: q = 8'h04;
            12'h1F4: q = 8'h04;
            12'h1F5: q = 8'h1F;
            12'h1F6: q = 8'h00;
            12'h1F7: q = 8'h00;
            12'h1F8: q = 8'h00;
            12'h1F9: q = 8'h00;
            12'h1FA: q = 8'h3E;
            12'h1FB: q = 8'h08;
            12'h1FC: q = 8'h08;
            12'h1FD: q = 8'h08;
            12'h1FE: q = 8'h08;
            12'h1FF: q = 8'h08;
            12'h200: q = 8'h08;
            12'h201: q = 8'h09;
            12'h202: q = 8'h07;
            12'h203: q = 8'h00;
            12'h204: q = 8'h00;
            12'h205: q = 8'h00;
            12'h206: q = 8'h37;
            12'h207: q = 8'h12;
            12'h208: q = 8'h0A;
            12'h209: q = 8'h06;
            12'h20A: q = 8'h0A;
            12'h20B: q = 8'h0A;
            12'h20C: q = 8'h12;
            12'h20D: q = 8'h37;
            12'h20E: q = 8'h00;
            12'h20F: q = 8'h00;
            12'h210: q = 8'h00;
            12'h211: q = 8'h00;
            12'h212: q = 8'h07;
            12'h213: q = 8'h02;
            12'h214: q = 8'h02;
            12'h215: q = 8'h02;
            12'h216: q = 8'h02;
            12'h217: q = 8'h02;
            12'h218: q = 8'h22;
            12'h219: q = 8'h3F;
            12'h21A: q = 8'h00;
            12'h21B: q = 8'h00;
            12'h21C: q = 8'h00;
            12'h21D: q = 8'h00;
            12'h21E: q = 8'h1B;
            12'h21F: q = 8'h1B;
            12'h220: q = 8'h1B;
            12'h221: q = 8'h1B;
            12'h222: q = 8'h15;
            12'h223: q = 8'h15;
            12'h224: q = 8'h15;
            12'h225: q = 8'h15;
            12'h226: q = 8'h00;
            12'h227: q = 8'h00;
            12'h228: q = 8'h00;
            12'h229: q = 8'h00;
            12'h22A: q = 8'h3B;
            12'h22B: q = 8'h12;
            12'h22C: q = 8'h16;
            12'h22D: q = 8'h16;
            12'h22E: q = 8'h1A;
            12'h22F: q = 8'h1A;
            12'h230: q = 8'h12;
            12'h231: q = 8'h17;
            12'h232: q = 8'h00;
            12'h233: q = 8'h00;
            12'h234: q = 8'h00;
            12'h235: q = 8'h00;
            12'h236: q = 8'h0E;
            12'h237: q = 8'h11;
            12'h238: q = 8'h11;
            12'h239: q = 8'h11;
            12'h23A: q = 8'h11;
            12'h23B: q = 8'h11;
            12'h23C: q = 8'h11;
            12'h23D: q = 8'h0E;
            12'h23E: q = 8'h00;
            12'h23F: q = 8'h00;
            12'h240: q = 8'h00;
            12'h241: q = 8'h00;
            12'h242: q = 8'h0F;
            12'h243: q = 8'h12;
            12'h244: q = 8'h12;
            12'h245: q = 8'h0E;
            12'h246: q = 8'h02;
            12'h247: q = 8'h02;
            12'h248: q = 8'h02;
            12'h249: q = 8'h07;
            12'h24A: q = 8'h00;
            12'h24B: q = 8'h00;
            12'h24C: q = 8'h00;
            12'h24D: q = 8'h00;
            12'h24E: q = 8'h0E;
            12'h24F: q = 8'h11;
            12'h250: q = 8'h11;
            12'h251: q = 8'h11;
            12'h252: q = 8'h11;
            12'h253: q = 8'h17;
            12'h254: q = 8'h19;
            12'h255: q = 8'h0E;
            12'h256: q = 8'h18;
            12'h257: q = 8'h00;
            12'h258: q = 8'h00;
            12'h259: q = 8'h00;
            12'h25A: q = 8'h0F;
            12'h25B: q = 8'h12;
            12'h25C: q = 8'h12;
            12'h25D: q = 8'h0E;
            12'h25E: q = 8'h0A;
            12'h25F: q = 8'h12;
            12'h260: q = 8'h12;
            12'h261: q = 8'h37;
            12'h262: q = 8'h00;
            12'h263: q = 8'h00;
            12'h264: q = 8'h00;
            12'h265: q = 8'h00;
            12'h266: q = 8'h1E;
            12'h267: q = 8'h11;
            12'h268: q = 8'h01;
            12'h269: q = 8'h06;
            12'h26A: q = 8'h08;
            12'h26B: q = 8'h10;
            12'h26C: q = 8'h11;
            12'h26D: q = 8'h0F;
            12'h26E: q = 8'h00;
            12'h26F: q = 8'h00;
            12'h270: q = 8'h00;
            12'h271: q = 8'h00;
            12'h272: q = 8'h1F;
            12'h273: q = 8'h15;
            12'h274: q = 8'h04;
            12'h275: q = 8'h04;
            12'h276: q = 8'h04;
            12'h277: q = 8'h04;
            12'h278: q = 8'h04;
            12'h279: q = 8'h0E;
            12'h27A: q = 8'h00;
            12'h27B: q = 8'h00;
            12'h27C: q = 8'h00;
            12'h27D: q = 8'h00;
            12'h27E: q = 8'h33;
            12'h27F: q = 8'h12;
            12'h280: q = 8'h12;
            12'h281: q = 8'h12;
            12'h282: q = 8'h12;
            12'h283: q = 8'h12;
            12'h284: q = 8'h12;
            12'h285: q = 8'h0C;
            12'h286: q = 8'h00;
            12'h287: q = 8'h00;
            12'h288: q = 8'h00;
            12'h289: q = 8'h00;
            12'h28A: q = 8'h33;
            12'h28B: q = 8'h12;
            12'h28C: q = 8'h12;
            12'h28D: q = 8'h0A;
            12'h28E: q = 8'h0A;
            12'h28F: q = 8'h0C;
            12'h290: q = 8'h04;
            12'h291: q = 8'h04;
            12'h292: q = 8'h00;
            12'h293: q = 8'h00;
            12'h294: q = 8'h00;
            12'h295: q = 8'h00;
            12'h296: q = 8'h15;
            12'h297: q = 8'h15;
            12'h298: q = 8'h15;
            12'h299: q = 8'h0E;
            12'h29A: q = 8'h0A;
            12'h29B: q = 8'h0A;
            12'h29C: q = 8'h0A;
            12'h29D: q = 8'h0A;
            12'h29E: q = 8'h00;
            12'h29F: q = 8'h00;
            12'h2A0: q = 8'h00;
            12'h2A1: q = 8'h00;
            12'h2A2: q = 8'h1B;
            12'h2A3: q = 8'h0A;
            12'h2A4: q = 8'h0A;
            12'h2A5: q = 8'h04;
            12'h2A6: q = 8'h04;
            12'h2A7: q = 8'h0A;
            12'h2A8: q = 8'h0A;
            12'h2A9: q = 8'h1B;
            12'h2AA: q = 8'h00;
            12'h2AB: q = 8'h00;
            12'h2AC: q = 8'h00;
            12'h2AD: q = 8'h00;
            12'h2AE: q = 8'h1B;
            12'h2AF: q = 8'h0A;
            12'h2B0: q = 8'h0A;
            12'h2B1: q = 8'h04;
            12'h2B2: q = 8'h04;
            12'h2B3: q = 8'h04;
            12'h2B4: q = 8'h04;
            12'h2B5: q = 8'h0E;
            12'h2B6: q = 8'h00;
            12'h2B7: q = 8'h00;
            12'h2B8: q = 8'h00;
            12'h2B9: q = 8'h00;
            12'h2BA: q = 8'h1F;
            12'h2BB: q = 8'h09;
            12'h2BC: q = 8'h08;
            12'h2BD: q = 8'h04;
            12'h2BE: q = 8'h04;
            12'h2BF: q = 8'h02;
            12'h2C0: q = 8'h12;
            12'h2C1: q = 8'h1F;
            12'h2C2: q = 8'h00;
            12'h2C3: q = 8'h00;
            12'h2C4: q = 8'h00;
            12'h2C5: q = 8'h1C;
            12'h2C6: q = 8'h04;
            12'h2C7: q = 8'h04;
            12'h2C8: q = 8'h04;
            12'h2C9: q = 8'h04;
            12'h2CA: q = 8'h04;
            12'h2CB: q = 8'h04;
            12'h2CC: q = 8'h04;
            12'h2CD: q = 8'h04;
            12'h2CE: q = 8'h1C;
            12'h2CF: q = 8'h00;
            12'h2D0: q = 8'h00;
            12'h2D1: q = 8'h02;
            12'h2D2: q = 8'h02;
            12'h2D3: q = 8'h02;
            12'h2D4: q = 8'h04;
            12'h2D5: q = 8'h04;
            12'h2D6: q = 8'h08;
            12'h2D7: q = 8'h08;
            12'h2D8: q = 8'h08;
            12'h2D9: q = 8'h10;
            12'h2DA: q = 8'h00;
            12'h2DB: q = 8'h00;
            12'h2DC: q = 8'h00;
            12'h2DD: q = 8'h0E;
            12'h2DE: q = 8'h08;
            12'h2DF: q = 8'h08;
            12'h2E0: q = 8'h08;
            12'h2E1: q = 8'h08;
            12'h2E2: q = 8'h08;
            12'h2E3: q = 8'h08;
            12'h2E4: q = 8'h08;
            12'h2E5: q = 8'h08;
            12'h2E6: q = 8'h0E;
            12'h2E7: q = 8'h00;
            12'h2E8: q = 8'h00;
            12'h2E9: q = 8'h04;
            12'h2EA: q = 8'h0A;
            12'h2EB: q = 8'h00;
            12'h2EC: q = 8'h00;
            12'h2ED: q = 8'h00;
            12'h2EE: q = 8'h00;
            12'h2EF: q = 8'h00;
            12'h2F0: q = 8'h00;
            12'h2F1: q = 8'h00;
            12'h2F2: q = 8'h00;
            12'h2F3: q = 8'h00;
            12'h2F4: q = 8'h00;
            12'h2F5: q = 8'h00;
            12'h2F6: q = 8'h00;
            12'h2F7: q = 8'h00;
            12'h2F8: q = 8'h00;
            12'h2F9: q = 8'h00;
            12'h2FA: q = 8'h00;
            12'h2FB: q = 8'h00;
            12'h2FC: q = 8'h00;
            12'h2FD: q = 8'h00;
            12'h2FE: q = 8'h00;
            12'h2FF: q = 8'h3F;
            12'h300: q = 8'h00;
            12'h301: q = 8'h04;
            12'h302: q = 8'h00;
            12'h303: q = 8'h00;
            12'h304: q = 8'h00;
            12'h305: q = 8'h00;
            12'h306: q = 8'h00;
            12'h307: q = 8'h00;
            12'h308: q = 8'h00;
            12'h309: q = 8'h00;
            12'h30A: q = 8'h00;
            12'h30B: q = 8'h00;
            12'h30C: q = 8'h00;
            12'h30D: q = 8'h00;
            12'h30E: q = 8'h00;
            12'h30F: q = 8'h00;
            12'h310: q = 8'h00;
            12'h311: q = 8'h0C;
            12'h312: q = 8'h12;
            12'h313: q = 8'h1C;
            12'h314: q = 8'h12;
            12'h315: q = 8'h3C;
            12'h316: q = 8'h00;
            12'h317: q = 8'h00;
            12'h318: q = 8'h00;
            12'h319: q = 8'h00;
            12'h31A: q = 8'h03;
            12'h31B: q = 8'h02;
            12'h31C: q = 8'h02;
            12'h31D: q = 8'h0E;
            12'h31E: q = 8'h12;
            12'h31F: q = 8'h12;
            12'h320: q = 8'h12;
            12'h321: q = 8'h0E;
            12'h322: q = 8'h00;
            12'h323: q = 8'h00;
            12'h324: q = 8'h00;
            12'h325: q = 8'h00;
            12'h326: q = 8'h00;
            12'h327: q = 8'h00;
            12'h328: q = 8'h00;
            12'h329: q = 8'h1C;
            12'h32A: q = 8'h12;
            12'h32B: q = 8'h02;
            12'h32C: q = 8'h02;
            12'h32D: q = 8'h1C;
            12'h32E: q = 8'h00;
            12'h32F: q = 8'h00;
            12'h330: q = 8'h00;
            12'h331: q = 8'h00;
            12'h332: q = 8'h18;
            12'h333: q = 8'h10;
            12'h334: q = 8'h10;
            12'h335: q = 8'h1C;
            12'h336: q = 8'h12;
            12'h337: q = 8'h12;
            12'h338: q = 8'h12;
            12'h339: q = 8'h3C;
            12'h33A: q = 8'h00;
            12'h33B: q = 8'h00;
            12'h33C: q = 8'h00;
            12'h33D: q = 8'h00;
            12'h33E: q = 8'h00;
            12'h33F: q = 8'h00;
            12'h340: q = 8'h00;
            12'h341: q = 8'h0C;
            12'h342: q = 8'h12;
            12'h343: q = 8'h1E;
            12'h344: q = 8'h02;
            12'h345: q = 8'h1C;
            12'h346: q = 8'h00;
            12'h347: q = 8'h00;
            12'h348: q = 8'h00;
            12'h349: q = 8'h00;
            12'h34A: q = 8'h38;
            12'h34B: q = 8'h04;
            12'h34C: q = 8'h04;
            12'h34D: q = 8'h1E;
            12'h34E: q = 8'h04;
            12'h34F: q = 8'h04;
            12'h350: q = 8'h04;
            12'h351: q = 8'h1E;
            12'h352: q = 8'h00;
            12'h353: q = 8'h00;
            12'h354: q = 8'h00;
            12'h355: q = 8'h00;
            12'h356: q = 8'h00;
            12'h357: q = 8'h00;
            12'h358: q = 8'h00;
            12'h359: q = 8'h3C;
            12'h35A: q = 8'h12;
            12'h35B: q = 8'h0C;
            12'h35C: q = 8'h02;
            12'h35D: q = 8'h1E;
            12'h35E: q = 8'h22;
            12'h35F: q = 8'h1C;
            12'h360: q = 8'h00;
            12'h361: q = 8'h00;
            12'h362: q = 8'h03;
            12'h363: q = 8'h02;
            12'h364: q = 8'h02;
            12'h365: q = 8'h0E;
            12'h366: q = 8'h12;
            12'h367: q = 8'h12;
            12'h368: q = 8'h12;
            12'h369: q = 8'h37;
            12'h36A: q = 8'h00;
            12'h36B: q = 8'h00;
            12'h36C: q = 8'h00;
            12'h36D: q = 8'h00;
            12'h36E: q = 8'h04;
            12'h36F: q = 8'h00;
            12'h370: q = 8'h00;
            12'h371: q = 8'h06;
            12'h372: q = 8'h04;
            12'h373: q = 8'h04;
            12'h374: q = 8'h04;
            12'h375: q = 8'h0E;
            12'h376: q = 8'h00;
            12'h377: q = 8'h00;
            12'h378: q = 8'h00;
            12'h379: q = 8'h00;
            12'h37A: q = 8'h08;
            12'h37B: q = 8'h00;
            12'h37C: q = 8'h00;
            12'h37D: q = 8'h0C;
            12'h37E: q = 8'h08;
            12'h37F: q = 8'h08;
            12'h380: q = 8'h08;
            12'h381: q = 8'h08;
            12'h382: q = 8'h08;
            12'h383: q = 8'h07;
            12'h384: q = 8'h00;
            12'h385: q = 8'h00;
            12'h386: q = 8'h03;
            12'h387: q = 8'h02;
            12'h388: q = 8'h02;
            12'h389: q = 8'h3A;
            12'h38A: q = 8'h0A;
            12'h38B: q = 8'h0E;
            12'h38C: q = 8'h12;
            12'h38D: q = 8'h37;
            12'h38E: q = 8'h00;
            12'h38F: q = 8'h00;
            12'h390: q = 8'h00;
            12'h391: q = 8'h00;
            12'h392: q = 8'h07;
            12'h393: q = 8'h04;
            12'h394: q = 8'h04;
            12'h395: q = 8'h04;
            12'h396: q = 8'h04;
            12'h397: q = 8'h04;
            12'h398: q = 8'h04;
            12'h399: q = 8'h1F;
            12'h39A: q = 8'h00;
            12'h39B: q = 8'h00;
            12'h39C: q = 8'h00;
            12'h39D: q = 8'h00;
            12'h39E: q = 8'h00;
            12'h39F: q = 8'h00;
            12'h3A0: q = 8'h00;
            12'h3A1: q = 8'h0F;
            12'h3A2: q = 8'h15;
            12'h3A3: q = 8'h15;
            12'h3A4: q = 8'h15;
            12'h3A5: q = 8'h15;
            12'h3A6: q = 8'h00;
            12'h3A7: q = 8'h00;
            12'h3A8: q = 8'h00;
            12'h3A9: q = 8'h00;
            12'h3AA: q = 8'h00;
            12'h3AB: q = 8'h00;
            12'h3AC: q = 8'h00;
            12'h3AD: q = 8'h0F;
            12'h3AE: q = 8'h12;
            12'h3AF: q = 8'h12;
            12'h3B0: q = 8'h12;
            12'h3B1: q = 8'h37;
            12'h3B2: q = 8'h00;
            12'h3B3: q = 8'h00;
            12'h3B4: q = 8'h00;
            12'h3B5: q = 8'h00;
            12'h3B6: q = 8'h00;
            12'h3B7: q = 8'h00;
            12'h3B8: q = 8'h00;
            12'h3B9: q = 8'h0C;
            12'h3BA: q = 8'h12;
            12'h3BB: q = 8'h12;
            12'h3BC: q = 8'h12;
            12'h3BD: q = 8'h0C;
            12'h3BE: q = 8'h00;
            12'h3BF: q = 8'h00;
            12'h3C0: q = 8'h00;
            12'h3C1: q = 8'h00;
            12'h3C2: q = 8'h00;
            12'h3C3: q = 8'h00;
            12'h3C4: q = 8'h00;
            12'h3C5: q = 8'h0F;
            12'h3C6: q = 8'h12;
            12'h3C7: q = 8'h12;
            12'h3C8: q = 8'h12;
            12'h3C9: q = 8'h0E;
            12'h3CA: q = 8'h02;
            12'h3CB: q = 8'h07;
            12'h3CC: q = 8'h00;
            12'h3CD: q = 8'h00;
            12'h3CE: q = 8'h00;
            12'h3CF: q = 8'h00;
            12'h3D0: q = 8'h00;
            12'h3D1: q = 8'h1C;
            12'h3D2: q = 8'h12;
            12'h3D3: q = 8'h12;
            12'h3D4: q = 8'h12;
            12'h3D5: q = 8'h1C;
            12'h3D6: q = 8'h10;
            12'h3D7: q = 8'h38;
            12'h3D8: q = 8'h00;
            12'h3D9: q = 8'h00;
            12'h3DA: q = 8'h00;
            12'h3DB: q = 8'h00;
            12'h3DC: q = 8'h00;
            12'h3DD: q = 8'h1B;
            12'h3DE: q = 8'h06;
            12'h3DF: q = 8'h02;
            12'h3E0: q = 8'h02;
            12'h3E1: q = 8'h07;
            12'h3E2: q = 8'h00;
            12'h3E3: q = 8'h00;
            12'h3E4: q = 8'h00;
            12'h3E5: q = 8'h00;
            12'h3E6: q = 8'h00;
            12'h3E7: q = 8'h00;
            12'h3E8: q = 8'h00;
            12'h3E9: q = 8'h1E;
            12'h3EA: q = 8'h02;
            12'h3EB: q = 8'h0C;
            12'h3EC: q = 8'h10;
            12'h3ED: q = 8'h1E;
            12'h3EE: q = 8'h00;
            12'h3EF: q = 8'h00;
            12'h3F0: q = 8'h00;
            12'h3F1: q = 8'h00;
            12'h3F2: q = 8'h00;
            12'h3F3: q = 8'h04;
            12'h3F4: q = 8'h04;
            12'h3F5: q = 8'h0E;
            12'h3F6: q = 8'h04;
            12'h3F7: q = 8'h04;
            12'h3F8: q = 8'h04;
            12'h3F9: q = 8'h18;
            12'h3FA: q = 8'h00;
            12'h3FB: q = 8'h00;
            12'h3FC: q = 8'h00;
            12'h3FD: q = 8'h00;
            12'h3FE: q = 8'h00;
            12'h3FF: q = 8'h00;
            12'h400: q = 8'h00;
            12'h401: q = 8'h1B;
            12'h402: q = 8'h12;
            12'h403: q = 8'h12;
            12'h404: q = 8'h12;
            12'h405: q = 8'h3C;
            12'h406: q = 8'h00;
            12'h407: q = 8'h00;
            12'h408: q = 8'h00;
            12'h409: q = 8'h00;
            12'h40A: q = 8'h00;
            12'h40B: q = 8'h00;
            12'h40C: q = 8'h00;
            12'h40D: q = 8'h37;
            12'h40E: q = 8'h12;
            12'h40F: q = 8'h0A;
            12'h410: q = 8'h0C;
            12'h411: q = 8'h04;
            12'h412: q = 8'h00;
            12'h413: q = 8'h00;
            12'h414: q = 8'h00;
            12'h415: q = 8'h00;
            12'h416: q = 8'h00;
            12'h417: q = 8'h00;
            12'h418: q = 8'h00;
            12'h419: q = 8'h15;
            12'h41A: q = 8'h15;
            12'h41B: q = 8'h0E;
            12'h41C: q = 8'h0A;
            12'h41D: q = 8'h0A;
            12'h41E: q = 8'h00;
            12'h41F: q = 8'h00;
            12'h420: q = 8'h00;
            12'h421: q = 8'h00;
            12'h422: q = 8'h00;
            12'h423: q = 8'h00;
            12'h424: q = 8'h00;
            12'h425: q = 8'h1B;
            12'h426: q = 8'h0A;
            12'h427: q = 8'h04;
            12'h428: q = 8'h0A;
            12'h429: q = 8'h1B;
            12'h42A: q = 8'h00;
            12'h42B: q = 8'h00;
            12'h42C: q = 8'h00;
            12'h42D: q = 8'h00;
            12'h42E: q = 8'h00;
            12'h42F: q = 8'h00;
            12'h430: q = 8'h00;
            12'h431: q = 8'h37;
            12'h432: q = 8'h12;
            12'h433: q = 8'h0A;
            12'h434: q = 8'h0C;
            12'h435: q = 8'h04;
            12'h436: q = 8'h04;
            12'h437: q = 8'h03;
            12'h438: q = 8'h00;
            12'h439: q = 8'h00;
            12'h43A: q = 8'h00;
            12'h43B: q = 8'h00;
            12'h43C: q = 8'h00;
            12'h43D: q = 8'h1E;
            12'h43E: q = 8'h08;
            12'h43F: q = 8'h04;
            12'h440: q = 8'h04;
            12'h441: q = 8'h1E;
            12'h442: q = 8'h00;
            12'h443: q = 8'h00;
            12'h444: q = 8'h00;
            12'h445: q = 8'h18;
            12'h446: q = 8'h08;
            12'h447: q = 8'h08;
            12'h448: q = 8'h08;
            12'h449: q = 8'h04;
            12'h44A: q = 8'h08;
            12'h44B: q = 8'h08;
            12'h44C: q = 8'h08;
            12'h44D: q = 8'h08;
            12'h44E: q = 8'h18;
            12'h44F: q = 8'h00;
            12'h450: q = 8'h08;
            12'h451: q = 8'h08;
            12'h452: q = 8'h08;
            12'h453: q = 8'h08;
            12'h454: q = 8'h08;
            12'h455: q = 8'h08;
            12'h456: q = 8'h08;
            12'h457: q = 8'h08;
            12'h458: q = 8'h08;
            12'h459: q = 8'h08;
            12'h45A: q = 8'h08;
            12'h45B: q = 8'h08;
            12'h45C: q = 8'h00;
            12'h45D: q = 8'h06;
            12'h45E: q = 8'h04;
            12'h45F: q = 8'h04;
            12'h460: q = 8'h04;
            12'h461: q = 8'h08;
            12'h462: q = 8'h04;
            12'h463: q = 8'h04;
            12'h464: q = 8'h04;
            12'h465: q = 8'h04;
            12'h466: q = 8'h06;
            12'h467: q = 8'h00;
            12'h468: q = 8'h02;
            12'h469: q = 8'h25;
            12'h46A: q = 8'h18;
            12'h46B: q = 8'h00;
            12'h46C: q = 8'h00;
            12'h46D: q = 8'h00;
            12'h46E: q = 8'h00;
            12'h46F: q = 8'h00;
            12'h470: q = 8'h00;
            12'h471: q = 8'h00;
            12'h472: q = 8'h00;
            12'h473: q = 8'h00;
            12'h474: q = 8'h00;
            12'h475: q = 8'h00;
            12'h476: q = 8'h00;
            12'h477: q = 8'h00;
            12'h478: q = 8'h00;
            12'h479: q = 8'h00;
            12'h47A: q = 8'h00;
            12'h47B: q = 8'h00;
            12'h47C: q = 8'h00;
            12'h47D: q = 8'h00;
            12'h47E: q = 8'h00;
            12'h47F: q = 8'h00;
            12'h480: q = 8'h00;
            12'h481: q = 8'h00;
            12'h482: q = 8'h00;
            12'h483: q = 8'h00;
            12'h484: q = 8'h00;
            12'h485: q = 8'h00;
            12'h486: q = 8'h00;
            12'h487: q = 8'h08;
            12'h488: q = 8'h08;
            12'h489: q = 8'h08;
            12'h48A: q = 8'h08;
            12'h48B: q = 8'h08;
            12'h48C: q = 8'h08;
            12'h48D: q = 8'h08;
            12'h48E: q = 8'h00;
            12'h48F: q = 8'h00;
            12'h490: q = 8'h18;
            12'h491: q = 8'h18;
            12'h492: q = 8'h00;
            12'h493: q = 8'h00;
            12'h494: q = 8'h00;
            12'h495: q = 8'h48;
            12'h496: q = 8'h6C;
            12'h497: q = 8'h24;
            12'h498: q = 8'h12;
            12'h499: q = 8'h00;
            12'h49A: q = 8'h00;
            12'h49B: q = 8'h00;
            12'h49C: q = 8'h00;
            12'h49D: q = 8'h00;
            12'h49E: q = 8'h00;
            12'h49F: q = 8'h00;
            12'h4A0: q = 8'h00;
            12'h4A1: q = 8'h00;
            12'h4A2: q = 8'h00;
            12'h4A3: q = 8'h00;
            12'h4A4: q = 8'h00;
            12'h4A5: q = 8'h00;
            12'h4A6: q = 8'h00;
            12'h4A7: q = 8'h24;
            12'h4A8: q = 8'h24;
            12'h4A9: q = 8'h24;
            12'h4AA: q = 8'h7F;
            12'h4AB: q = 8'h12;
            12'h4AC: q = 8'h12;
            12'h4AD: q = 8'h12;
            12'h4AE: q = 8'h7F;
            12'h4AF: q = 8'h12;
            12'h4B0: q = 8'h12;
            12'h4B1: q = 8'h12;
            12'h4B2: q = 8'h00;
            12'h4B3: q = 8'h00;
            12'h4B4: q = 8'h00;
            12'h4B5: q = 8'h00;
            12'h4B6: q = 8'h08;
            12'h4B7: q = 8'h1C;
            12'h4B8: q = 8'h2A;
            12'h4B9: q = 8'h2A;
            12'h4BA: q = 8'h0A;
            12'h4BB: q = 8'h0C;
            12'h4BC: q = 8'h18;
            12'h4BD: q = 8'h28;
            12'h4BE: q = 8'h28;
            12'h4BF: q = 8'h2A;
            12'h4C0: q = 8'h2A;
            12'h4C1: q = 8'h1C;
            12'h4C2: q = 8'h08;
            12'h4C3: q = 8'h08;
            12'h4C4: q = 8'h00;
            12'h4C5: q = 8'h00;
            12'h4C6: q = 8'h00;
            12'h4C7: q = 8'h22;
            12'h4C8: q = 8'h25;
            12'h4C9: q = 8'h15;
            12'h4CA: q = 8'h15;
            12'h4CB: q = 8'h15;
            12'h4CC: q = 8'h2A;
            12'h4CD: q = 8'h58;
            12'h4CE: q = 8'h54;
            12'h4CF: q = 8'h54;
            12'h4D0: q = 8'h54;
            12'h4D1: q = 8'h22;
            12'h4D2: q = 8'h00;
            12'h4D3: q = 8'h00;
            12'h4D4: q = 8'h00;
            12'h4D5: q = 8'h00;
            12'h4D6: q = 8'h00;
            12'h4D7: q = 8'h0C;
            12'h4D8: q = 8'h12;
            12'h4D9: q = 8'h12;
            12'h4DA: q = 8'h12;
            12'h4DB: q = 8'h0A;
            12'h4DC: q = 8'h76;
            12'h4DD: q = 8'h25;
            12'h4DE: q = 8'h29;
            12'h4DF: q = 8'h11;
            12'h4E0: q = 8'h91;
            12'h4E1: q = 8'h6E;
            12'h4E2: q = 8'h00;
            12'h4E3: q = 8'h00;
            12'h4E4: q = 8'h00;
            12'h4E5: q = 8'h06;
            12'h4E6: q = 8'h06;
            12'h4E7: q = 8'h04;
            12'h4E8: q = 8'h03;
            12'h4E9: q = 8'h00;
            12'h4EA: q = 8'h00;
            12'h4EB: q = 8'h00;
            12'h4EC: q = 8'h00;
            12'h4ED: q = 8'h00;
            12'h4EE: q = 8'h00;
            12'h4EF: q = 8'h00;
            12'h4F0: q = 8'h00;
            12'h4F1: q = 8'h00;
            12'h4F2: q = 8'h00;
            12'h4F3: q = 8'h00;
            12'h4F4: q = 8'h00;
            12'h4F5: q = 8'h40;
            12'h4F6: q = 8'h20;
            12'h4F7: q = 8'h10;
            12'h4F8: q = 8'h10;
            12'h4F9: q = 8'h08;
            12'h4FA: q = 8'h08;
            12'h4FB: q = 8'h08;
            12'h4FC: q = 8'h08;
            12'h4FD: q = 8'h08;
            12'h4FE: q = 8'h08;
            12'h4FF: q = 8'h10;
            12'h500: q = 8'h10;
            12'h501: q = 8'h20;
            12'h502: q = 8'h40;
            12'h503: q = 8'h00;
            12'h504: q = 8'h00;
            12'h505: q = 8'h02;
            12'h506: q = 8'h04;
            12'h507: q = 8'h08;
            12'h508: q = 8'h08;
            12'h509: q = 8'h10;
            12'h50A: q = 8'h10;
            12'h50B: q = 8'h10;
            12'h50C: q = 8'h10;
            12'h50D: q = 8'h10;
            12'h50E: q = 8'h10;
            12'h50F: q = 8'h08;
            12'h510: q = 8'h08;
            12'h511: q = 8'h04;
            12'h512: q = 8'h02;
            12'h513: q = 8'h00;
            12'h514: q = 8'h00;
            12'h515: q = 8'h00;
            12'h516: q = 8'h00;
            12'h517: q = 8'h00;
            12'h518: q = 8'h08;
            12'h519: q = 8'h08;
            12'h51A: q = 8'h6B;
            12'h51B: q = 8'h1C;
            12'h51C: q = 8'h1C;
            12'h51D: q = 8'h6B;
            12'h51E: q = 8'h08;
            12'h51F: q = 8'h08;
            12'h520: q = 8'h00;
            12'h521: q = 8'h00;
            12'h522: q = 8'h00;
            12'h523: q = 8'h00;
            12'h524: q = 8'h00;
            12'h525: q = 8'h00;
            12'h526: q = 8'h00;
            12'h527: q = 8'h00;
            12'h528: q = 8'h08;
            12'h529: q = 8'h08;
            12'h52A: q = 8'h08;
            12'h52B: q = 8'h08;
            12'h52C: q = 8'h7F;
            12'h52D: q = 8'h08;
            12'h52E: q = 8'h08;
            12'h52F: q = 8'h08;
            12'h530: q = 8'h08;
            12'h531: q = 8'h00;
            12'h532: q = 8'h00;
            12'h533: q = 8'h00;
            12'h534: q = 8'h00;
            12'h535: q = 8'h00;
            12'h536: q = 8'h00;
            12'h537: q = 8'h00;
            12'h538: q = 8'h00;
            12'h539: q = 8'h00;
            12'h53A: q = 8'h00;
            12'h53B: q = 8'h00;
            12'h53C: q = 8'h00;
            12'h53D: q = 8'h00;
            12'h53E: q = 8'h00;
            12'h53F: q = 8'h00;
            12'h540: q = 8'h06;
            12'h541: q = 8'h06;
            12'h542: q = 8'h04;
            12'h543: q = 8'h03;
            12'h544: q = 8'h00;
            12'h545: q = 8'h00;
            12'h546: q = 8'h00;
            12'h547: q = 8'h00;
            12'h548: q = 8'h00;
            12'h549: q = 8'h00;
            12'h54A: q = 8'h00;
            12'h54B: q = 8'h00;
            12'h54C: q = 8'hFE;
            12'h54D: q = 8'h00;
            12'h54E: q = 8'h00;
            12'h54F: q = 8'h00;
            12'h550: q = 8'h00;
            12'h551: q = 8'h00;
            12'h552: q = 8'h00;
            12'h553: q = 8'h00;
            12'h554: q = 8'h00;
            12'h555: q = 8'h00;
            12'h556: q = 8'h00;
            12'h557: q = 8'h00;
            12'h558: q = 8'h00;
            12'h559: q = 8'h00;
            12'h55A: q = 8'h00;
            12'h55B: q = 8'h00;
            12'h55C: q = 8'h00;
            12'h55D: q = 8'h00;
            12'h55E: q = 8'h00;
            12'h55F: q = 8'h00;
            12'h560: q = 8'h06;
            12'h561: q = 8'h06;
            12'h562: q = 8'h00;
            12'h563: q = 8'h00;
            12'h564: q = 8'h00;
            12'h565: q = 8'h00;
            12'h566: q = 8'h80;
            12'h567: q = 8'h40;
            12'h568: q = 8'h40;
            12'h569: q = 8'h20;
            12'h56A: q = 8'h20;
            12'h56B: q = 8'h10;
            12'h56C: q = 8'h10;
            12'h56D: q = 8'h08;
            12'h56E: q = 8'h08;
            12'h56F: q = 8'h04;
            12'h570: q = 8'h04;
            12'h571: q = 8'h02;
            12'h572: q = 8'h02;
            12'h573: q = 8'h00;
            12'h574: q = 8'h00;
            12'h575: q = 8'h00;
            12'h576: q = 8'h00;
            12'h577: q = 8'h18;
            12'h578: q = 8'h24;
            12'h579: q = 8'h42;
            12'h57A: q = 8'h42;
            12'h57B: q = 8'h42;
            12'h57C: q = 8'h42;
            12'h57D: q = 8'h42;
            12'h57E: q = 8'h42;
            12'h57F: q = 8'h42;
            12'h580: q = 8'h24;
            12'h581: q = 8'h18;
            12'h582: q = 8'h00;
            12'h583: q = 8'h00;
            12'h584: q = 8'h00;
            12'h585: q = 8'h00;
            12'h586: q = 8'h00;
            12'h587: q = 8'h08;
            12'h588: q = 8'h0E;
            12'h589: q = 8'h08;
            12'h58A: q = 8'h08;
            12'h58B: q = 8'h08;
            12'h58C: q = 8'h08;
            12'h58D: q = 8'h08;
            12'h58E: q = 8'h08;
            12'h58F: q = 8'h08;
            12'h590: q = 8'h08;
            12'h591: q = 8'h3E;
            12'h592: q = 8'h00;
            12'h593: q = 8'h00;
            12'h594: q = 8'h00;
            12'h595: q = 8'h00;
            12'h596: q = 8'h00;
            12'h597: q = 8'h3C;
            12'h598: q = 8'h42;
            12'h599: q = 8'h42;
            12'h59A: q = 8'h42;
            12'h59B: q = 8'h20;
            12'h59C: q = 8'h20;
            12'h59D: q = 8'h10;
            12'h59E: q = 8'h08;
            12'h59F: q = 8'h04;
            12'h5A0: q = 8'h42;
            12'h5A1: q = 8'h7E;
            12'h5A2: q = 8'h00;
            12'h5A3: q = 8'h00;
            12'h5A4: q = 8'h00;
            12'h5A5: q = 8'h00;
            12'h5A6: q = 8'h00;
            12'h5A7: q = 8'h3C;
            12'h5A8: q = 8'h42;
            12'h5A9: q = 8'h42;
            12'h5AA: q = 8'h20;
            12'h5AB: q = 8'h18;
            12'h5AC: q = 8'h20;
            12'h5AD: q = 8'h40;
            12'h5AE: q = 8'h40;
            12'h5AF: q = 8'h42;
            12'h5B0: q = 8'h22;
            12'h5B1: q = 8'h1C;
            12'h5B2: q = 8'h00;
            12'h5B3: q = 8'h00;
            12'h5B4: q = 8'h00;
            12'h5B5: q = 8'h00;
            12'h5B6: q = 8'h00;
            12'h5B7: q = 8'h20;
            12'h5B8: q = 8'h30;
            12'h5B9: q = 8'h28;
            12'h5BA: q = 8'h24;
            12'h5BB: q = 8'h24;
            12'h5BC: q = 8'h22;
            12'h5BD: q = 8'h22;
            12'h5BE: q = 8'h7E;
            12'h5BF: q = 8'h20;
            12'h5C0: q = 8'h20;
            12'h5C1: q = 8'h78;
            12'h5C2: q = 8'h00;
            12'h5C3: q = 8'h00;
            12'h5C4: q = 8'h00;
            12'h5C5: q = 8'h00;
            12'h5C6: q = 8'h00;
            12'h5C7: q = 8'h7E;
            12'h5C8: q = 8'h02;
            12'h5C9: q = 8'h02;
            12'h5CA: q = 8'h02;
            12'h5CB: q = 8'h1A;
            12'h5CC: q = 8'h26;
            12'h5CD: q = 8'h40;
            12'h5CE: q = 8'h40;
            12'h5CF: q = 8'h42;
            12'h5D0: q = 8'h22;
            12'h5D1: q = 8'h1C;
            12'h5D2: q = 8'h00;
            12'h5D3: q = 8'h00;
            12'h5D4: q = 8'h00;
            12'h5D5: q = 8'h00;
            12'h5D6: q = 8'h00;
            12'h5D7: q = 8'h38;
            12'h5D8: q = 8'h24;
            12'h5D9: q = 8'h02;
            12'h5DA: q = 8'h02;
            12'h5DB: q = 8'h1A;
            12'h5DC: q = 8'h26;
            12'h5DD: q = 8'h42;
            12'h5DE: q = 8'h42;
            12'h5DF: q = 8'h42;
            12'h5E0: q = 8'h24;
            12'h5E1: q = 8'h18;
            12'h5E2: q = 8'h00;
            12'h5E3: q = 8'h00;
            12'h5E4: q = 8'h00;
            12'h5E5: q = 8'h00;
            12'h5E6: q = 8'h00;
            12'h5E7: q = 8'h7E;
            12'h5E8: q = 8'h22;
            12'h5E9: q = 8'h22;
            12'h5EA: q = 8'h10;
            12'h5EB: q = 8'h10;
            12'h5EC: q = 8'h08;
            12'h5ED: q = 8'h08;
            12'h5EE: q = 8'h08;
            12'h5EF: q = 8'h08;
            12'h5F0: q = 8'h08;
            12'h5F1: q = 8'h08;
            12'h5F2: q = 8'h00;
            12'h5F3: q = 8'h00;
            12'h5F4: q = 8'h00;
            12'h5F5: q = 8'h00;
            12'h5F6: q = 8'h00;
            12'h5F7: q = 8'h3C;
            12'h5F8: q = 8'h42;
            12'h5F9: q = 8'h42;
            12'h5FA: q = 8'h42;
            12'h5FB: q = 8'h24;
            12'h5FC: q = 8'h18;
            12'h5FD: q = 8'h24;
            12'h5FE: q = 8'h42;
            12'h5FF: q = 8'h42;
            12'h600: q = 8'h42;
            12'h601: q = 8'h3C;
            12'h602: q = 8'h00;
            12'h603: q = 8'h00;
            12'h604: q = 8'h00;
            12'h605: q = 8'h00;
            12'h606: q = 8'h00;
            12'h607: q = 8'h18;
            12'h608: q = 8'h24;
            12'h609: q = 8'h42;
            12'h60A: q = 8'h42;
            12'h60B: q = 8'h42;
            12'h60C: q = 8'h64;
            12'h60D: q = 8'h58;
            12'h60E: q = 8'h40;
            12'h60F: q = 8'h40;
            12'h610: q = 8'h24;
            12'h611: q = 8'h1C;
            12'h612: q = 8'h00;
            12'h613: q = 8'h00;
            12'h614: q = 8'h00;
            12'h615: q = 8'h00;
            12'h616: q = 8'h00;
            12'h617: q = 8'h00;
            12'h618: q = 8'h00;
            12'h619: q = 8'h00;
            12'h61A: q = 8'h18;
            12'h61B: q = 8'h18;
            12'h61C: q = 8'h00;
            12'h61D: q = 8'h00;
            12'h61E: q = 8'h00;
            12'h61F: q = 8'h00;
            12'h620: q = 8'h18;
            12'h621: q = 8'h18;
            12'h622: q = 8'h00;
            12'h623: q = 8'h00;
            12'h624: q = 8'h00;
            12'h625: q = 8'h00;
            12'h626: q = 8'h00;
            12'h627: q = 8'h00;
            12'h628: q = 8'h00;
            12'h629: q = 8'h00;
            12'h62A: q = 8'h00;
            12'h62B: q = 8'h08;
            12'h62C: q = 8'h00;
            12'h62D: q = 8'h00;
            12'h62E: q = 8'h00;
            12'h62F: q = 8'h00;
            12'h630: q = 8'h00;
            12'h631: q = 8'h08;
            12'h632: q = 8'h08;
            12'h633: q = 8'h04;
            12'h634: q = 8'h00;
            12'h635: q = 8'h00;
            12'h636: q = 8'h00;
            12'h637: q = 8'h40;
            12'h638: q = 8'h20;
            12'h639: q = 8'h10;
            12'h63A: q = 8'h08;
            12'h63B: q = 8'h04;
            12'h63C: q = 8'h02;
            12'h63D: q = 8'h04;
            12'h63E: q = 8'h08;
            12'h63F: q = 8'h10;
            12'h640: q = 8'h20;
            12'h641: q = 8'h40;
            12'h642: q = 8'h00;
            12'h643: q = 8'h00;
            12'h644: q = 8'h00;
            12'h645: q = 8'h00;
            12'h646: q = 8'h00;
            12'h647: q = 8'h00;
            12'h648: q = 8'h00;
            12'h649: q = 8'h00;
            12'h64A: q = 8'h7F;
            12'h64B: q = 8'h00;
            12'h64C: q = 8'h00;
            12'h64D: q = 8'h00;
            12'h64E: q = 8'h7F;
            12'h64F: q = 8'h00;
            12'h650: q = 8'h00;
            12'h651: q = 8'h00;
            12'h652: q = 8'h00;
            12'h653: q = 8'h00;
            12'h654: q = 8'h00;
            12'h655: q = 8'h00;
            12'h656: q = 8'h00;
            12'h657: q = 8'h02;
            12'h658: q = 8'h04;
            12'h659: q = 8'h08;
            12'h65A: q = 8'h10;
            12'h65B: q = 8'h20;
            12'h65C: q = 8'h40;
            12'h65D: q = 8'h20;
            12'h65E: q = 8'h10;
            12'h65F: q = 8'h08;
            12'h660: q = 8'h04;
            12'h661: q = 8'h02;
            12'h662: q = 8'h00;
            12'h663: q = 8'h00;
            12'h664: q = 8'h00;
            12'h665: q = 8'h00;
            12'h666: q = 8'h00;
            12'h667: q = 8'h3C;
            12'h668: q = 8'h42;
            12'h669: q = 8'h42;
            12'h66A: q = 8'h46;
            12'h66B: q = 8'h40;
            12'h66C: q = 8'h20;
            12'h66D: q = 8'h10;
            12'h66E: q = 8'h10;
            12'h66F: q = 8'h00;
            12'h670: q = 8'h18;
            12'h671: q = 8'h18;
            12'h672: q = 8'h00;
            12'h673: q = 8'h00;
            12'h674: q = 8'h00;
            12'h675: q = 8'h00;
            12'h676: q = 8'h00;
            12'h677: q = 8'h1C;
            12'h678: q = 8'h22;
            12'h679: q = 8'h5A;
            12'h67A: q = 8'h55;
            12'h67B: q = 8'h55;
            12'h67C: q = 8'h55;
            12'h67D: q = 8'h55;
            12'h67E: q = 8'h2D;
            12'h67F: q = 8'h42;
            12'h680: q = 8'h22;
            12'h681: q = 8'h1C;
            12'h682: q = 8'h00;
            12'h683: q = 8'h00;
            12'h684: q = 8'h00;
            12'h685: q = 8'h00;
            12'h686: q = 8'h00;
            12'h687: q = 8'h08;
            12'h688: q = 8'h08;
            12'h689: q = 8'h18;
            12'h68A: q = 8'h14;
            12'h68B: q = 8'h14;
            12'h68C: q = 8'h24;
            12'h68D: q = 8'h3C;
            12'h68E: q = 8'h22;
            12'h68F: q = 8'h42;
            12'h690: q = 8'h42;
            12'h691: q = 8'hE7;
            12'h692: q = 8'h00;
            12'h693: q = 8'h00;
            12'h694: q = 8'h00;
            12'h695: q = 8'h00;
            12'h696: q = 8'h00;
            12'h697: q = 8'h1F;
            12'h698: q = 8'h22;
            12'h699: q = 8'h22;
            12'h69A: q = 8'h22;
            12'h69B: q = 8'h1E;
            12'h69C: q = 8'h22;
            12'h69D: q = 8'h42;
            12'h69E: q = 8'h42;
            12'h69F: q = 8'h42;
            12'h6A0: q = 8'h22;
            12'h6A1: q = 8'h1F;
            12'h6A2: q = 8'h00;
            12'h6A3: q = 8'h00;
            12'h6A4: q = 8'h00;
            12'h6A5: q = 8'h00;
            12'h6A6: q = 8'h00;
            12'h6A7: q = 8'h7C;
            12'h6A8: q = 8'h42;
            12'h6A9: q = 8'h42;
            12'h6AA: q = 8'h01;
            12'h6AB: q = 8'h01;
            12'h6AC: q = 8'h01;
            12'h6AD: q = 8'h01;
            12'h6AE: q = 8'h01;
            12'h6AF: q = 8'h42;
            12'h6B0: q = 8'h22;
            12'h6B1: q = 8'h1C;
            12'h6B2: q = 8'h00;
            12'h6B3: q = 8'h00;
            12'h6B4: q = 8'h00;
            12'h6B5: q = 8'h00;
            12'h6B6: q = 8'h00;
            12'h6B7: q = 8'h1F;
            12'h6B8: q = 8'h22;
            12'h6B9: q = 8'h42;
            12'h6BA: q = 8'h42;
            12'h6BB: q = 8'h42;
            12'h6BC: q = 8'h42;
            12'h6BD: q = 8'h42;
            12'h6BE: q = 8'h42;
            12'h6BF: q = 8'h42;
            12'h6C0: q = 8'h22;
            12'h6C1: q = 8'h1F;
            12'h6C2: q = 8'h00;
            12'h6C3: q = 8'h00;
            12'h6C4: q = 8'h00;
            12'h6C5: q = 8'h00;
            12'h6C6: q = 8'h00;
            12'h6C7: q = 8'h3F;
            12'h6C8: q = 8'h42;
            12'h6C9: q = 8'h12;
            12'h6CA: q = 8'h12;
            12'h6CB: q = 8'h1E;
            12'h6CC: q = 8'h12;
            12'h6CD: q = 8'h12;
            12'h6CE: q = 8'h02;
            12'h6CF: q = 8'h42;
            12'h6D0: q = 8'h42;
            12'h6D1: q = 8'h3F;
            12'h6D2: q = 8'h00;
            12'h6D3: q = 8'h00;
            12'h6D4: q = 8'h00;
            12'h6D5: q = 8'h00;
            12'h6D6: q = 8'h00;
            12'h6D7: q = 8'h3F;
            12'h6D8: q = 8'h42;
            12'h6D9: q = 8'h12;
            12'h6DA: q = 8'h12;
            12'h6DB: q = 8'h1E;
            12'h6DC: q = 8'h12;
            12'h6DD: q = 8'h12;
            12'h6DE: q = 8'h02;
            12'h6DF: q = 8'h02;
            12'h6E0: q = 8'h02;
            12'h6E1: q = 8'h07;
            12'h6E2: q = 8'h00;
            12'h6E3: q = 8'h00;
            12'h6E4: q = 8'h00;
            12'h6E5: q = 8'h00;
            12'h6E6: q = 8'h00;
            12'h6E7: q = 8'h3C;
            12'h6E8: q = 8'h22;
            12'h6E9: q = 8'h22;
            12'h6EA: q = 8'h01;
            12'h6EB: q = 8'h01;
            12'h6EC: q = 8'h01;
            12'h6ED: q = 8'h71;
            12'h6EE: q = 8'h21;
            12'h6EF: q = 8'h22;
            12'h6F0: q = 8'h22;
            12'h6F1: q = 8'h1C;
            12'h6F2: q = 8'h00;
            12'h6F3: q = 8'h00;
            12'h6F4: q = 8'h00;
            12'h6F5: q = 8'h00;
            12'h6F6: q = 8'h00;
            12'h6F7: q = 8'hE7;
            12'h6F8: q = 8'h42;
            12'h6F9: q = 8'h42;
            12'h6FA: q = 8'h42;
            12'h6FB: q = 8'h42;
            12'h6FC: q = 8'h7E;
            12'h6FD: q = 8'h42;
            12'h6FE: q = 8'h42;
            12'h6FF: q = 8'h42;
            12'h700: q = 8'h42;
            12'h701: q = 8'hE7;
            12'h702: q = 8'h00;
            12'h703: q = 8'h00;
            12'h704: q = 8'h00;
            12'h705: q = 8'h00;
            12'h706: q = 8'h00;
            12'h707: q = 8'h3E;
            12'h708: q = 8'h08;
            12'h709: q = 8'h08;
            12'h70A: q = 8'h08;
            12'h70B: q = 8'h08;
            12'h70C: q = 8'h08;
            12'h70D: q = 8'h08;
            12'h70E: q = 8'h08;
            12'h70F: q = 8'h08;
            12'h710: q = 8'h08;
            12'h711: q = 8'h3E;
            12'h712: q = 8'h00;
            12'h713: q = 8'h00;
            12'h714: q = 8'h00;
            12'h715: q = 8'h00;
            12'h716: q = 8'h00;
            12'h717: q = 8'h7C;
            12'h718: q = 8'h10;
            12'h719: q = 8'h10;
            12'h71A: q = 8'h10;
            12'h71B: q = 8'h10;
            12'h71C: q = 8'h10;
            12'h71D: q = 8'h10;
            12'h71E: q = 8'h10;
            12'h71F: q = 8'h10;
            12'h720: q = 8'h10;
            12'h721: q = 8'h10;
            12'h722: q = 8'h11;
            12'h723: q = 8'h0F;
            12'h724: q = 8'h00;
            12'h725: q = 8'h00;
            12'h726: q = 8'h00;
            12'h727: q = 8'h77;
            12'h728: q = 8'h22;
            12'h729: q = 8'h12;
            12'h72A: q = 8'h0A;
            12'h72B: q = 8'h0E;
            12'h72C: q = 8'h0A;
            12'h72D: q = 8'h12;
            12'h72E: q = 8'h12;
            12'h72F: q = 8'h22;
            12'h730: q = 8'h22;
            12'h731: q = 8'h77;
            12'h732: q = 8'h00;
            12'h733: q = 8'h00;
            12'h734: q = 8'h00;
            12'h735: q = 8'h00;
            12'h736: q = 8'h00;
            12'h737: q = 8'h07;
            12'h738: q = 8'h02;
            12'h739: q = 8'h02;
            12'h73A: q = 8'h02;
            12'h73B: q = 8'h02;
            12'h73C: q = 8'h02;
            12'h73D: q = 8'h02;
            12'h73E: q = 8'h02;
            12'h73F: q = 8'h02;
            12'h740: q = 8'h42;
            12'h741: q = 8'h7F;
            12'h742: q = 8'h00;
            12'h743: q = 8'h00;
            12'h744: q = 8'h00;
            12'h745: q = 8'h00;
            12'h746: q = 8'h00;
            12'h747: q = 8'h77;
            12'h748: q = 8'h36;
            12'h749: q = 8'h36;
            12'h74A: q = 8'h36;
            12'h74B: q = 8'h36;
            12'h74C: q = 8'h2A;
            12'h74D: q = 8'h2A;
            12'h74E: q = 8'h2A;
            12'h74F: q = 8'h2A;
            12'h750: q = 8'h2A;
            12'h751: q = 8'h6B;
            12'h752: q = 8'h00;
            12'h753: q = 8'h00;
            12'h754: q = 8'h00;
            12'h755: q = 8'h00;
            12'h756: q = 8'h00;
            12'h757: q = 8'hE3;
            12'h758: q = 8'h46;
            12'h759: q = 8'h46;
            12'h75A: q = 8'h4A;
            12'h75B: q = 8'h4A;
            12'h75C: q = 8'h52;
            12'h75D: q = 8'h52;
            12'h75E: q = 8'h52;
            12'h75F: q = 8'h62;
            12'h760: q = 8'h62;
            12'h761: q = 8'h47;
            12'h762: q = 8'h00;
            12'h763: q = 8'h00;
            12'h764: q = 8'h00;
            12'h765: q = 8'h00;
            12'h766: q = 8'h00;
            12'h767: q = 8'h1C;
            12'h768: q = 8'h22;
            12'h769: q = 8'h41;
            12'h76A: q = 8'h41;
            12'h76B: q = 8'h41;
            12'h76C: q = 8'h41;
            12'h76D: q = 8'h41;
            12'h76E: q = 8'h41;
            12'h76F: q = 8'h41;
            12'h770: q = 8'h22;
            12'h771: q = 8'h1C;
            12'h772: q = 8'h00;
            12'h773: q = 8'h00;
            12'h774: q = 8'h00;
            12'h775: q = 8'h00;
            12'h776: q = 8'h00;
            12'h777: q = 8'h3F;
            12'h778: q = 8'h42;
            12'h779: q = 8'h42;
            12'h77A: q = 8'h42;
            12'h77B: q = 8'h42;
            12'h77C: q = 8'h3E;
            12'h77D: q = 8'h02;
            12'h77E: q = 8'h02;
            12'h77F: q = 8'h02;
            12'h780: q = 8'h02;
            12'h781: q = 8'h07;
            12'h782: q = 8'h00;
            12'h783: q = 8'h00;
            12'h784: q = 8'h00;
            12'h785: q = 8'h00;
            12'h786: q = 8'h00;
            12'h787: q = 8'h1C;
            12'h788: q = 8'h22;
            12'h789: q = 8'h41;
            12'h78A: q = 8'h41;
            12'h78B: q = 8'h41;
            12'h78C: q = 8'h41;
            12'h78D: q = 8'h41;
            12'h78E: q = 8'h4D;
            12'h78F: q = 8'h53;
            12'h790: q = 8'h32;
            12'h791: q = 8'h1C;
            12'h792: q = 8'h60;
            12'h793: q = 8'h00;
            12'h794: q = 8'h00;
            12'h795: q = 8'h00;
            12'h796: q = 8'h00;
            12'h797: q = 8'h3F;
            12'h798: q = 8'h42;
            12'h799: q = 8'h42;
            12'h79A: q = 8'h42;
            12'h79B: q = 8'h3E;
            12'h79C: q = 8'h12;
            12'h79D: q = 8'h12;
            12'h79E: q = 8'h22;
            12'h79F: q = 8'h22;
            12'h7A0: q = 8'h42;
            12'h7A1: q = 8'hC7;
            12'h7A2: q = 8'h00;
            12'h7A3: q = 8'h00;
            12'h7A4: q = 8'h00;
            12'h7A5: q = 8'h00;
            12'h7A6: q = 8'h00;
            12'h7A7: q = 8'h7C;
            12'h7A8: q = 8'h42;
            12'h7A9: q = 8'h42;
            12'h7AA: q = 8'h02;
            12'h7AB: q = 8'h04;
            12'h7AC: q = 8'h18;
            12'h7AD: q = 8'h20;
            12'h7AE: q = 8'h40;
            12'h7AF: q = 8'h42;
            12'h7B0: q = 8'h42;
            12'h7B1: q = 8'h3E;
            12'h7B2: q = 8'h00;
            12'h7B3: q = 8'h00;
            12'h7B4: q = 8'h00;
            12'h7B5: q = 8'h00;
            12'h7B6: q = 8'h00;
            12'h7B7: q = 8'h7F;
            12'h7B8: q = 8'h49;
            12'h7B9: q = 8'h08;
            12'h7BA: q = 8'h08;
            12'h7BB: q = 8'h08;
            12'h7BC: q = 8'h08;
            12'h7BD: q = 8'h08;
            12'h7BE: q = 8'h08;
            12'h7BF: q = 8'h08;
            12'h7C0: q = 8'h08;
            12'h7C1: q = 8'h1C;
            12'h7C2: q = 8'h00;
            12'h7C3: q = 8'h00;
            12'h7C4: q = 8'h00;
            12'h7C5: q = 8'h00;
            12'h7C6: q = 8'h00;
            12'h7C7: q = 8'hE7;
            12'h7C8: q = 8'h42;
            12'h7C9: q = 8'h42;
            12'h7CA: q = 8'h42;
            12'h7CB: q = 8'h42;
            12'h7CC: q = 8'h42;
            12'h7CD: q = 8'h42;
            12'h7CE: q = 8'h42;
            12'h7CF: q = 8'h42;
            12'h7D0: q = 8'h42;
            12'h7D1: q = 8'h3C;
            12'h7D2: q = 8'h00;
            12'h7D3: q = 8'h00;
            12'h7D4: q = 8'h00;
            12'h7D5: q = 8'h00;
            12'h7D6: q = 8'h00;
            12'h7D7: q = 8'hE7;
            12'h7D8: q = 8'h42;
            12'h7D9: q = 8'h42;
            12'h7DA: q = 8'h22;
            12'h7DB: q = 8'h24;
            12'h7DC: q = 8'h24;
            12'h7DD: q = 8'h14;
            12'h7DE: q = 8'h14;
            12'h7DF: q = 8'h18;
            12'h7E0: q = 8'h08;
            12'h7E1: q = 8'h08;
            12'h7E2: q = 8'h00;
            12'h7E3: q = 8'h00;
            12'h7E4: q = 8'h00;
            12'h7E5: q = 8'h00;
            12'h7E6: q = 8'h00;
            12'h7E7: q = 8'h6B;
            12'h7E8: q = 8'h49;
            12'h7E9: q = 8'h49;
            12'h7EA: q = 8'h49;
            12'h7EB: q = 8'h49;
            12'h7EC: q = 8'h55;
            12'h7ED: q = 8'h55;
            12'h7EE: q = 8'h36;
            12'h7EF: q = 8'h22;
            12'h7F0: q = 8'h22;
            12'h7F1: q = 8'h22;
            12'h7F2: q = 8'h00;
            12'h7F3: q = 8'h00;
            12'h7F4: q = 8'h00;
            12'h7F5: q = 8'h00;
            12'h7F6: q = 8'h00;
            12'h7F7: q = 8'hE7;
            12'h7F8: q = 8'h42;
            12'h7F9: q = 8'h24;
            12'h7FA: q = 8'h24;
            12'h7FB: q = 8'h18;
            12'h7FC: q = 8'h18;
            12'h7FD: q = 8'h18;
            12'h7FE: q = 8'h24;
            12'h7FF: q = 8'h24;
            12'h800: q = 8'h42;
            12'h801: q = 8'hE7;
            12'h802: q = 8'h00;
            12'h803: q = 8'h00;
            12'h804: q = 8'h00;
            12'h805: q = 8'h00;
            12'h806: q = 8'h00;
            12'h807: q = 8'h77;
            12'h808: q = 8'h22;
            12'h809: q = 8'h22;
            12'h80A: q = 8'h14;
            12'h80B: q = 8'h14;
            12'h80C: q = 8'h08;
            12'h80D: q = 8'h08;
            12'h80E: q = 8'h08;
            12'h80F: q = 8'h08;
            12'h810: q = 8'h08;
            12'h811: q = 8'h1C;
            12'h812: q = 8'h00;
            12'h813: q = 8'h00;
            12'h814: q = 8'h00;
            12'h815: q = 8'h00;
            12'h816: q = 8'h00;
            12'h817: q = 8'h7E;
            12'h818: q = 8'h21;
            12'h819: q = 8'h20;
            12'h81A: q = 8'h10;
            12'h81B: q = 8'h10;
            12'h81C: q = 8'h08;
            12'h81D: q = 8'h04;
            12'h81E: q = 8'h04;
            12'h81F: q = 8'h42;
            12'h820: q = 8'h42;
            12'h821: q = 8'h3F;
            12'h822: q = 8'h00;
            12'h823: q = 8'h00;
            12'h824: q = 8'h00;
            12'h825: q = 8'h78;
            12'h826: q = 8'h08;
            12'h827: q = 8'h08;
            12'h828: q = 8'h08;
            12'h829: q = 8'h08;
            12'h82A: q = 8'h08;
            12'h82B: q = 8'h08;
            12'h82C: q = 8'h08;
            12'h82D: q = 8'h08;
            12'h82E: q = 8'h08;
            12'h82F: q = 8'h08;
            12'h830: q = 8'h08;
            12'h831: q = 8'h08;
            12'h832: q = 8'h78;
            12'h833: q = 8'h00;
            12'h834: q = 8'h00;
            12'h835: q = 8'h00;
            12'h836: q = 8'h02;
            12'h837: q = 8'h02;
            12'h838: q = 8'h04;
            12'h839: q = 8'h04;
            12'h83A: q = 8'h08;
            12'h83B: q = 8'h08;
            12'h83C: q = 8'h08;
            12'h83D: q = 8'h10;
            12'h83E: q = 8'h10;
            12'h83F: q = 8'h20;
            12'h840: q = 8'h20;
            12'h841: q = 8'h20;
            12'h842: q = 8'h40;
            12'h843: q = 8'h40;
            12'h844: q = 8'h00;
            12'h845: q = 8'h1E;
            12'h846: q = 8'h10;
            12'h847: q = 8'h10;
            12'h848: q = 8'h10;
            12'h849: q = 8'h10;
            12'h84A: q = 8'h10;
            12'h84B: q = 8'h10;
            12'h84C: q = 8'h10;
            12'h84D: q = 8'h10;
            12'h84E: q = 8'h10;
            12'h84F: q = 8'h10;
            12'h850: q = 8'h10;
            12'h851: q = 8'h10;
            12'h852: q = 8'h1E;
            12'h853: q = 8'h00;
            12'h854: q = 8'h00;
            12'h855: q = 8'h38;
            12'h856: q = 8'h44;
            12'h857: q = 8'h00;
            12'h858: q = 8'h00;
            12'h859: q = 8'h00;
            12'h85A: q = 8'h00;
            12'h85B: q = 8'h00;
            12'h85C: q = 8'h00;
            12'h85D: q = 8'h00;
            12'h85E: q = 8'h00;
            12'h85F: q = 8'h00;
            12'h860: q = 8'h00;
            12'h861: q = 8'h00;
            12'h862: q = 8'h00;
            12'h863: q = 8'h00;
            12'h864: q = 8'h00;
            12'h865: q = 8'h00;
            12'h866: q = 8'h00;
            12'h867: q = 8'h00;
            12'h868: q = 8'h00;
            12'h869: q = 8'h00;
            12'h86A: q = 8'h00;
            12'h86B: q = 8'h00;
            12'h86C: q = 8'h00;
            12'h86D: q = 8'h00;
            12'h86E: q = 8'h00;
            12'h86F: q = 8'h00;
            12'h870: q = 8'h00;
            12'h871: q = 8'h00;
            12'h872: q = 8'h00;
            12'h873: q = 8'hFF;
            12'h874: q = 8'h00;
            12'h875: q = 8'h06;
            12'h876: q = 8'h08;
            12'h877: q = 8'h00;
            12'h878: q = 8'h00;
            12'h879: q = 8'h00;
            12'h87A: q = 8'h00;
            12'h87B: q = 8'h00;
            12'h87C: q = 8'h00;
            12'h87D: q = 8'h00;
            12'h87E: q = 8'h00;
            12'h87F: q = 8'h00;
            12'h880: q = 8'h00;
            12'h881: q = 8'h00;
            12'h882: q = 8'h00;
            12'h883: q = 8'h00;
            12'h884: q = 8'h00;
            12'h885: q = 8'h00;
            12'h886: q = 8'h00;
            12'h887: q = 8'h00;
            12'h888: q = 8'h00;
            12'h889: q = 8'h00;
            12'h88A: q = 8'h00;
            12'h88B: q = 8'h3C;
            12'h88C: q = 8'h42;
            12'h88D: q = 8'h78;
            12'h88E: q = 8'h44;
            12'h88F: q = 8'h42;
            12'h890: q = 8'h42;
            12'h891: q = 8'hFC;
            12'h892: q = 8'h00;
            12'h893: q = 8'h00;
            12'h894: q = 8'h00;
            12'h895: q = 8'h00;
            12'h896: q = 8'h00;
            12'h897: q = 8'h03;
            12'h898: q = 8'h02;
            12'h899: q = 8'h02;
            12'h89A: q = 8'h02;
            12'h89B: q = 8'h1A;
            12'h89C: q = 8'h26;
            12'h89D: q = 8'h42;
            12'h89E: q = 8'h42;
            12'h89F: q = 8'h42;
            12'h8A0: q = 8'h26;
            12'h8A1: q = 8'h1A;
            12'h8A2: q = 8'h00;
            12'h8A3: q = 8'h00;
            12'h8A4: q = 8'h00;
            12'h8A5: q = 8'h00;
            12'h8A6: q = 8'h00;
            12'h8A7: q = 8'h00;
            12'h8A8: q = 8'h00;
            12'h8A9: q = 8'h00;
            12'h8AA: q = 8'h00;
            12'h8AB: q = 8'h38;
            12'h8AC: q = 8'h44;
            12'h8AD: q = 8'h02;
            12'h8AE: q = 8'h02;
            12'h8AF: q = 8'h02;
            12'h8B0: q = 8'h44;
            12'h8B1: q = 8'h38;
            12'h8B2: q = 8'h00;
            12'h8B3: q = 8'h00;
            12'h8B4: q = 8'h00;
            12'h8B5: q = 8'h00;
            12'h8B6: q = 8'h00;
            12'h8B7: q = 8'h60;
            12'h8B8: q = 8'h40;
            12'h8B9: q = 8'h40;
            12'h8BA: q = 8'h40;
            12'h8BB: q = 8'h78;
            12'h8BC: q = 8'h44;
            12'h8BD: q = 8'h42;
            12'h8BE: q = 8'h42;
            12'h8BF: q = 8'h42;
            12'h8C0: q = 8'h64;
            12'h8C1: q = 8'hD8;
            12'h8C2: q = 8'h00;
            12'h8C3: q = 8'h00;
            12'h8C4: q = 8'h00;
            12'h8C5: q = 8'h00;
            12'h8C6: q = 8'h00;
            12'h8C7: q = 8'h00;
            12'h8C8: q = 8'h00;
            12'h8C9: q = 8'h00;
            12'h8CA: q = 8'h00;
            12'h8CB: q = 8'h3C;
            12'h8CC: q = 8'h42;
            12'h8CD: q = 8'h7E;
            12'h8CE: q = 8'h02;
            12'h8CF: q = 8'h02;
            12'h8D0: q = 8'h42;
            12'h8D1: q = 8'h3C;
            12'h8D2: q = 8'h00;
            12'h8D3: q = 8'h00;
            12'h8D4: q = 8'h00;
            12'h8D5: q = 8'h00;
            12'h8D6: q = 8'h00;
            12'h8D7: q = 8'hF0;
            12'h8D8: q = 8'h88;
            12'h8D9: q = 8'h08;
            12'h8DA: q = 8'h08;
            12'h8DB: q = 8'h7E;
            12'h8DC: q = 8'h08;
            12'h8DD: q = 8'h08;
            12'h8DE: q = 8'h08;
            12'h8DF: q = 8'h08;
            12'h8E0: q = 8'h08;
            12'h8E1: q = 8'h3E;
            12'h8E2: q = 8'h00;
            12'h8E3: q = 8'h00;
            12'h8E4: q = 8'h00;
            12'h8E5: q = 8'h00;
            12'h8E6: q = 8'h00;
            12'h8E7: q = 8'h00;
            12'h8E8: q = 8'h00;
            12'h8E9: q = 8'h00;
            12'h8EA: q = 8'h00;
            12'h8EB: q = 8'h7C;
            12'h8EC: q = 8'h22;
            12'h8ED: q = 8'h22;
            12'h8EE: q = 8'h1C;
            12'h8EF: q = 8'h02;
            12'h8F0: q = 8'h3C;
            12'h8F1: q = 8'h42;
            12'h8F2: q = 8'h42;
            12'h8F3: q = 8'h3C;
            12'h8F4: q = 8'h00;
            12'h8F5: q = 8'h00;
            12'h8F6: q = 8'h00;
            12'h8F7: q = 8'h03;
            12'h8F8: q = 8'h02;
            12'h8F9: q = 8'h02;
            12'h8FA: q = 8'h02;
            12'h8FB: q = 8'h3A;
            12'h8FC: q = 8'h46;
            12'h8FD: q = 8'h42;
            12'h8FE: q = 8'h42;
            12'h8FF: q = 8'h42;
            12'h900: q = 8'h42;
            12'h901: q = 8'hE7;
            12'h902: q = 8'h00;
            12'h903: q = 8'h00;
            12'h904: q = 8'h00;
            12'h905: q = 8'h00;
            12'h906: q = 8'h00;
            12'h907: q = 8'h0C;
            12'h908: q = 8'h0C;
            12'h909: q = 8'h00;
            12'h90A: q = 8'h00;
            12'h90B: q = 8'h0E;
            12'h90C: q = 8'h08;
            12'h90D: q = 8'h08;
            12'h90E: q = 8'h08;
            12'h90F: q = 8'h08;
            12'h910: q = 8'h08;
            12'h911: q = 8'h3E;
            12'h912: q = 8'h00;
            12'h913: q = 8'h00;
            12'h914: q = 8'h00;
            12'h915: q = 8'h00;
            12'h916: q = 8'h00;
            12'h917: q = 8'h30;
            12'h918: q = 8'h30;
            12'h919: q = 8'h00;
            12'h91A: q = 8'h00;
            12'h91B: q = 8'h38;
            12'h91C: q = 8'h20;
            12'h91D: q = 8'h20;
            12'h91E: q = 8'h20;
            12'h91F: q = 8'h20;
            12'h920: q = 8'h20;
            12'h921: q = 8'h20;
            12'h922: q = 8'h22;
            12'h923: q = 8'h1E;
            12'h924: q = 8'h00;
            12'h925: q = 8'h00;
            12'h926: q = 8'h00;
            12'h927: q = 8'h03;
            12'h928: q = 8'h02;
            12'h929: q = 8'h02;
            12'h92A: q = 8'h02;
            12'h92B: q = 8'h72;
            12'h92C: q = 8'h12;
            12'h92D: q = 8'h0A;
            12'h92E: q = 8'h16;
            12'h92F: q = 8'h12;
            12'h930: q = 8'h22;
            12'h931: q = 8'h77;
            12'h932: q = 8'h00;
            12'h933: q = 8'h00;
            12'h934: q = 8'h00;
            12'h935: q = 8'h00;
            12'h936: q = 8'h00;
            12'h937: q = 8'h0E;
            12'h938: q = 8'h08;
            12'h939: q = 8'h08;
            12'h93A: q = 8'h08;
            12'h93B: q = 8'h08;
            12'h93C: q = 8'h08;
            12'h93D: q = 8'h08;
            12'h93E: q = 8'h08;
            12'h93F: q = 8'h08;
            12'h940: q = 8'h08;
            12'h941: q = 8'h3E;
            12'h942: q = 8'h00;
            12'h943: q = 8'h00;
            12'h944: q = 8'h00;
            12'h945: q = 8'h00;
            12'h946: q = 8'h00;
            12'h947: q = 8'h00;
            12'h948: q = 8'h00;
            12'h949: q = 8'h00;
            12'h94A: q = 8'h00;
            12'h94B: q = 8'h7F;
            12'h94C: q = 8'h92;
            12'h94D: q = 8'h92;
            12'h94E: q = 8'h92;
            12'h94F: q = 8'h92;
            12'h950: q = 8'h92;
            12'h951: q = 8'hB7;
            12'h952: q = 8'h00;
            12'h953: q = 8'h00;
            12'h954: q = 8'h00;
            12'h955: q = 8'h00;
            12'h956: q = 8'h00;
            12'h957: q = 8'h00;
            12'h958: q = 8'h00;
            12'h959: q = 8'h00;
            12'h95A: q = 8'h00;
            12'h95B: q = 8'h3B;
            12'h95C: q = 8'h46;
            12'h95D: q = 8'h42;
            12'h95E: q = 8'h42;
            12'h95F: q = 8'h42;
            12'h960: q = 8'h42;
            12'h961: q = 8'hE7;
            12'h962: q = 8'h00;
            12'h963: q = 8'h00;
            12'h964: q = 8'h00;
            12'h965: q = 8'h00;
            12'h966: q = 8'h00;
            12'h967: q = 8'h00;
            12'h968: q = 8'h00;
            12'h969: q = 8'h00;
            12'h96A: q = 8'h00;
            12'h96B: q = 8'h3C;
            12'h96C: q = 8'h42;
            12'h96D: q = 8'h42;
            12'h96E: q = 8'h42;
            12'h96F: q = 8'h42;
            12'h970: q = 8'h42;
            12'h971: q = 8'h3C;
            12'h972: q = 8'h00;
            12'h973: q = 8'h00;
            12'h974: q = 8'h00;
            12'h975: q = 8'h00;
            12'h976: q = 8'h00;
            12'h977: q = 8'h00;
            12'h978: q = 8'h00;
            12'h979: q = 8'h00;
            12'h97A: q = 8'h00;
            12'h97B: q = 8'h1B;
            12'h97C: q = 8'h26;
            12'h97D: q = 8'h42;
            12'h97E: q = 8'h42;
            12'h97F: q = 8'h42;
            12'h980: q = 8'h22;
            12'h981: q = 8'h1E;
            12'h982: q = 8'h02;
            12'h983: q = 8'h07;
            12'h984: q = 8'h00;
            12'h985: q = 8'h00;
            12'h986: q = 8'h00;
            12'h987: q = 8'h00;
            12'h988: q = 8'h00;
            12'h989: q = 8'h00;
            12'h98A: q = 8'h00;
            12'h98B: q = 8'h78;
            12'h98C: q = 8'h44;
            12'h98D: q = 8'h42;
            12'h98E: q = 8'h42;
            12'h98F: q = 8'h42;
            12'h990: q = 8'h44;
            12'h991: q = 8'h78;
            12'h992: q = 8'h40;
            12'h993: q = 8'hE0;
            12'h994: q = 8'h00;
            12'h995: q = 8'h00;
            12'h996: q = 8'h00;
            12'h997: q = 8'h00;
            12'h998: q = 8'h00;
            12'h999: q = 8'h00;
            12'h99A: q = 8'h00;
            12'h99B: q = 8'h77;
            12'h99C: q = 8'h4C;
            12'h99D: q = 8'h04;
            12'h99E: q = 8'h04;
            12'h99F: q = 8'h04;
            12'h9A0: q = 8'h04;
            12'h9A1: q = 8'h1F;
            12'h9A2: q = 8'h00;
            12'h9A3: q = 8'h00;
            12'h9A4: q = 8'h00;
            12'h9A5: q = 8'h00;
            12'h9A6: q = 8'h00;
            12'h9A7: q = 8'h00;
            12'h9A8: q = 8'h00;
            12'h9A9: q = 8'h00;
            12'h9AA: q = 8'h00;
            12'h9AB: q = 8'h7C;
            12'h9AC: q = 8'h42;
            12'h9AD: q = 8'h02;
            12'h9AE: q = 8'h3C;
            12'h9AF: q = 8'h40;
            12'h9B0: q = 8'h42;
            12'h9B1: q = 8'h3E;
            12'h9B2: q = 8'h00;
            12'h9B3: q = 8'h00;
            12'h9B4: q = 8'h00;
            12'h9B5: q = 8'h00;
            12'h9B6: q = 8'h00;
            12'h9B7: q = 8'h00;
            12'h9B8: q = 8'h00;
            12'h9B9: q = 8'h08;
            12'h9BA: q = 8'h08;
            12'h9BB: q = 8'h3E;
            12'h9BC: q = 8'h08;
            12'h9BD: q = 8'h08;
            12'h9BE: q = 8'h08;
            12'h9BF: q = 8'h08;
            12'h9C0: q = 8'h08;
            12'h9C1: q = 8'h30;
            12'h9C2: q = 8'h00;
            12'h9C3: q = 8'h00;
            12'h9C4: q = 8'h00;
            12'h9C5: q = 8'h00;
            12'h9C6: q = 8'h00;
            12'h9C7: q = 8'h00;
            12'h9C8: q = 8'h00;
            12'h9C9: q = 8'h00;
            12'h9CA: q = 8'h00;
            12'h9CB: q = 8'h63;
            12'h9CC: q = 8'h42;
            12'h9CD: q = 8'h42;
            12'h9CE: q = 8'h42;
            12'h9CF: q = 8'h42;
            12'h9D0: q = 8'h62;
            12'h9D1: q = 8'hDC;
            12'h9D2: q = 8'h00;
            12'h9D3: q = 8'h00;
            12'h9D4: q = 8'h00;
            12'h9D5: q = 8'h00;
            12'h9D6: q = 8'h00;
            12'h9D7: q = 8'h00;
            12'h9D8: q = 8'h00;
            12'h9D9: q = 8'h00;
            12'h9DA: q = 8'h00;
            12'h9DB: q = 8'hE7;
            12'h9DC: q = 8'h42;
            12'h9DD: q = 8'h24;
            12'h9DE: q = 8'h24;
            12'h9DF: q = 8'h14;
            12'h9E0: q = 8'h08;
            12'h9E1: q = 8'h08;
            12'h9E2: q = 8'h00;
            12'h9E3: q = 8'h00;
            12'h9E4: q = 8'h00;
            12'h9E5: q = 8'h00;
            12'h9E6: q = 8'h00;
            12'h9E7: q = 8'h00;
            12'h9E8: q = 8'h00;
            12'h9E9: q = 8'h00;
            12'h9EA: q = 8'h00;
            12'h9EB: q = 8'hEB;
            12'h9EC: q = 8'h49;
            12'h9ED: q = 8'h49;
            12'h9EE: q = 8'h55;
            12'h9EF: q = 8'h55;
            12'h9F0: q = 8'h22;
            12'h9F1: q = 8'h22;
            12'h9F2: q = 8'h00;
            12'h9F3: q = 8'h00;
            12'h9F4: q = 8'h00;
            12'h9F5: q = 8'h00;
            12'h9F6: q = 8'h00;
            12'h9F7: q = 8'h00;
            12'h9F8: q = 8'h00;
            12'h9F9: q = 8'h00;
            12'h9FA: q = 8'h00;
            12'h9FB: q = 8'h76;
            12'h9FC: q = 8'h24;
            12'h9FD: q = 8'h18;
            12'h9FE: q = 8'h18;
            12'h9FF: q = 8'h18;
            12'hA00: q = 8'h24;
            12'hA01: q = 8'h6E;
            12'hA02: q = 8'h00;
            12'hA03: q = 8'h00;
            12'hA04: q = 8'h00;
            12'hA05: q = 8'h00;
            12'hA06: q = 8'h00;
            12'hA07: q = 8'h00;
            12'hA08: q = 8'h00;
            12'hA09: q = 8'h00;
            12'hA0A: q = 8'h00;
            12'hA0B: q = 8'hE7;
            12'hA0C: q = 8'h42;
            12'hA0D: q = 8'h24;
            12'hA0E: q = 8'h24;
            12'hA0F: q = 8'h14;
            12'hA10: q = 8'h18;
            12'hA11: q = 8'h08;
            12'hA12: q = 8'h08;
            12'hA13: q = 8'h07;
            12'hA14: q = 8'h00;
            12'hA15: q = 8'h00;
            12'hA16: q = 8'h00;
            12'hA17: q = 8'h00;
            12'hA18: q = 8'h00;
            12'hA19: q = 8'h00;
            12'hA1A: q = 8'h00;
            12'hA1B: q = 8'h7E;
            12'hA1C: q = 8'h22;
            12'hA1D: q = 8'h10;
            12'hA1E: q = 8'h08;
            12'hA1F: q = 8'h08;
            12'hA20: q = 8'h44;
            12'hA21: q = 8'h7E;
            12'hA22: q = 8'h00;
            12'hA23: q = 8'h00;
            12'hA24: q = 8'h00;
            12'hA25: q = 8'hC0;
            12'hA26: q = 8'h20;
            12'hA27: q = 8'h20;
            12'hA28: q = 8'h20;
            12'hA29: q = 8'h20;
            12'hA2A: q = 8'h20;
            12'hA2B: q = 8'h10;
            12'hA2C: q = 8'h20;
            12'hA2D: q = 8'h20;
            12'hA2E: q = 8'h20;
            12'hA2F: q = 8'h20;
            12'hA30: q = 8'h20;
            12'hA31: q = 8'h20;
            12'hA32: q = 8'hC0;
            12'hA33: q = 8'h00;
            12'hA34: q = 8'h10;
            12'hA35: q = 8'h10;
            12'hA36: q = 8'h10;
            12'hA37: q = 8'h10;
            12'hA38: q = 8'h10;
            12'hA39: q = 8'h10;
            12'hA3A: q = 8'h10;
            12'hA3B: q = 8'h10;
            12'hA3C: q = 8'h10;
            12'hA3D: q = 8'h10;
            12'hA3E: q = 8'h10;
            12'hA3F: q = 8'h10;
            12'hA40: q = 8'h10;
            12'hA41: q = 8'h10;
            12'hA42: q = 8'h10;
            12'hA43: q = 8'h10;
            12'hA44: q = 8'h00;
            12'hA45: q = 8'h06;
            12'hA46: q = 8'h08;
            12'hA47: q = 8'h08;
            12'hA48: q = 8'h08;
            12'hA49: q = 8'h08;
            12'hA4A: q = 8'h08;
            12'hA4B: q = 8'h10;
            12'hA4C: q = 8'h08;
            12'hA4D: q = 8'h08;
            12'hA4E: q = 8'h08;
            12'hA4F: q = 8'h08;
            12'hA50: q = 8'h08;
            12'hA51: q = 8'h08;
            12'hA52: q = 8'h06;
            12'hA53: q = 8'h00;
            12'hA54: q = 8'h0C;
            12'hA55: q = 8'h32;
            12'hA56: q = 8'hC2;
            12'hA57: q = 8'h00;
            12'hA58: q = 8'h00;
            12'hA59: q = 8'h00;
            12'hA5A: q = 8'h00;
            12'hA5B: q = 8'h00;
            12'hA5C: q = 8'h00;
            12'hA5D: q = 8'h00;
            12'hA5E: q = 8'h00;
            12'hA5F: q = 8'h00;
            12'hA60: q = 8'h00;
            12'hA61: q = 8'h00;
            12'hA62: q = 8'h00;
            12'hA63: q = 8'h00;
            12'hA64: q = 8'h00;
            12'hA65: q = 8'h00;
            12'hA66: q = 8'h00;
            12'hA67: q = 8'h00;
            12'hA68: q = 8'h00;
            12'hA69: q = 8'h00;
            12'hA6A: q = 8'h00;
            12'hA6B: q = 8'h00;
            12'hA6C: q = 8'h00;
            12'hA6D: q = 8'h00;
            12'hA6E: q = 8'h00;
            12'hA6F: q = 8'h00;
            12'hA70: q = 8'h00;
            12'hA71: q = 8'h00;
            12'hA72: q = 8'h00;
            12'hA73: q = 8'h00;
            12'hA74: q = 8'h00;
            12'hA75: q = 8'h00;
            12'hA76: q = 8'h00;
            12'hA77: q = 8'h00;
            12'hA78: q = 8'h00;
            12'hA79: q = 8'h00;
            12'hA7A: q = 8'h00;
            12'hA7B: q = 8'h00;
            12'hA7C: q = 8'h00;
            12'hA7D: q = 8'h00;
            12'hA7E: q = 8'h00;
            12'hA7F: q = 8'h00;
            12'hA80: q = 8'h00;
            12'hA81: q = 8'h00;
            12'hA82: q = 8'h00;
            12'hA83: q = 8'h00;
            12'hA84: q = 8'h00;
            12'hA85: q = 8'h00;
            12'hA86: q = 8'h00;
            12'hA87: q = 8'h00;
            12'hA88: q = 8'h00;
            12'hA89: q = 8'h00;
            12'hA8A: q = 8'h00;
            12'hA8B: q = 8'h00;
            12'hA8C: q = 8'h00;
            12'hA8D: q = 8'h00;
            12'hA8E: q = 8'h00;
            12'hA8F: q = 8'h00;
            12'hA90: q = 8'h00;
            12'hA91: q = 8'h00;
            12'hA92: q = 8'h00;
            12'hA93: q = 8'h00;
            12'hA94: q = 8'h00;
            12'hA95: q = 8'h00;
            12'hA96: q = 8'h00;
            12'hA97: q = 8'h00;
            12'hA98: q = 8'h00;
            12'hA99: q = 8'h00;
            12'hA9A: q = 8'h00;
            12'hA9B: q = 8'h00;
            12'hA9C: q = 8'h00;
            12'hA9D: q = 8'h00;
            12'hA9E: q = 8'h00;
            12'hA9F: q = 8'h00;
            12'hAA0: q = 8'h00;
            12'hAA1: q = 8'h00;
            12'hAA2: q = 8'h00;
            12'hAA3: q = 8'h00;
            12'hAA4: q = 8'h00;
            12'hAA5: q = 8'h00;
            12'hAA6: q = 8'h00;
            12'hAA7: q = 8'h00;
            12'hAA8: q = 8'h00;
            12'hAA9: q = 8'h00;
            12'hAAA: q = 8'h00;
            12'hAAB: q = 8'h00;
            12'hAAC: q = 8'h00;
            12'hAAD: q = 8'h00;
            12'hAAE: q = 8'h00;
            12'hAAF: q = 8'h00;
            12'hAB0: q = 8'h00;
            12'hAB1: q = 8'h00;
            12'hAB2: q = 8'h00;
            12'hAB3: q = 8'h00;
            12'hAB4: q = 8'h00;
            12'hAB5: q = 8'h00;
            12'hAB6: q = 8'h00;
            12'hAB7: q = 8'h00;
            12'hAB8: q = 8'h00;
            12'hAB9: q = 8'h00;
            12'hABA: q = 8'h00;
            12'hABB: q = 8'h00;
            12'hABC: q = 8'h00;
            12'hABD: q = 8'h00;
            12'hABE: q = 8'h00;
            12'hABF: q = 8'h00;
            12'hAC0: q = 8'h00;
            12'hAC1: q = 8'h00;
            12'hAC2: q = 8'h00;
            12'hAC3: q = 8'h00;
            12'hAC4: q = 8'h00;
            12'hAC5: q = 8'h00;
            12'hAC6: q = 8'h00;
            12'hAC7: q = 8'h00;
            12'hAC8: q = 8'h00;
            12'hAC9: q = 8'h00;
            12'hACA: q = 8'h00;
            12'hACB: q = 8'h00;
            12'hACC: q = 8'h00;
            12'hACD: q = 8'h00;
            12'hACE: q = 8'h00;
            12'hACF: q = 8'h00;
            12'hAD0: q = 8'h00;
            12'hAD1: q = 8'h00;
            12'hAD2: q = 8'h00;
            12'hAD3: q = 8'h00;
            12'hAD4: q = 8'h00;
            12'hAD5: q = 8'h00;
            12'hAD6: q = 8'h00;
            12'hAD7: q = 8'h00;
            12'hAD8: q = 8'h00;
            12'hAD9: q = 8'h00;
            12'hADA: q = 8'h00;
            12'hADB: q = 8'h00;
            12'hADC: q = 8'h00;
            12'hADD: q = 8'h00;
            12'hADE: q = 8'h00;
            12'hADF: q = 8'h00;
            12'hAE0: q = 8'h00;
            12'hAE1: q = 8'h00;
            12'hAE2: q = 8'h00;
            12'hAE3: q = 8'h00;
            12'hAE4: q = 8'h00;
            12'hAE5: q = 8'h00;
            12'hAE6: q = 8'h00;
            12'hAE7: q = 8'h00;
            12'hAE8: q = 8'h00;
            12'hAE9: q = 8'h00;
            12'hAEA: q = 8'h00;
            12'hAEB: q = 8'h00;
            12'hAEC: q = 8'h00;
            12'hAED: q = 8'h00;
            12'hAEE: q = 8'h00;
            12'hAEF: q = 8'h00;
            12'hAF0: q = 8'h00;
            12'hAF1: q = 8'h00;
            12'hAF2: q = 8'h00;
            12'hAF3: q = 8'h00;
            12'hAF4: q = 8'h00;
            12'hAF5: q = 8'h00;
            12'hAF6: q = 8'h00;
            12'hAF7: q = 8'h00;
            12'hAF8: q = 8'h00;
            12'hAF9: q = 8'h00;
            12'hAFA: q = 8'h00;
            12'hAFB: q = 8'h00;
            12'hAFC: q = 8'h00;
            12'hAFD: q = 8'h00;
            12'hAFE: q = 8'h00;
            12'hAFF: q = 8'h00;
            12'hB00: q = 8'h00;
            12'hB01: q = 8'h00;
            12'hB02: q = 8'h00;
            12'hB03: q = 8'h00;
            12'hB04: q = 8'h00;
            12'hB05: q = 8'h00;
            12'hB06: q = 8'h00;
            12'hB07: q = 8'h00;
            12'hB08: q = 8'h00;
            12'hB09: q = 8'h00;
            12'hB0A: q = 8'h00;
            12'hB0B: q = 8'h00;
            12'hB0C: q = 8'h00;
            12'hB0D: q = 8'h00;
            12'hB0E: q = 8'h00;
            12'hB0F: q = 8'h00;
            12'hB10: q = 8'h00;
            12'hB11: q = 8'h00;
            12'hB12: q = 8'h00;
            12'hB13: q = 8'h00;
            12'hB14: q = 8'h00;
            12'hB15: q = 8'h00;
            12'hB16: q = 8'h00;
            12'hB17: q = 8'h00;
            12'hB18: q = 8'h00;
            12'hB19: q = 8'h00;
            12'hB1A: q = 8'h00;
            12'hB1B: q = 8'h00;
            12'hB1C: q = 8'h00;
            12'hB1D: q = 8'h00;
            12'hB1E: q = 8'h00;
            12'hB1F: q = 8'h00;
            12'hB20: q = 8'h00;
            12'hB21: q = 8'h00;
            12'hB22: q = 8'h00;
            12'hB23: q = 8'h00;
            12'hB24: q = 8'h00;
            12'hB25: q = 8'h00;
            12'hB26: q = 8'h00;
            12'hB27: q = 8'h00;
            12'hB28: q = 8'h00;
            12'hB29: q = 8'h00;
            12'hB2A: q = 8'h00;
            12'hB2B: q = 8'h00;
            12'hB2C: q = 8'h00;
            12'hB2D: q = 8'h00;
            12'hB2E: q = 8'h00;
            12'hB2F: q = 8'h00;
            12'hB30: q = 8'h00;
            12'hB31: q = 8'h00;
            12'hB32: q = 8'h00;
            12'hB33: q = 8'h00;
            12'hB34: q = 8'h00;
            12'hB35: q = 8'h00;
            12'hB36: q = 8'h00;
            12'hB37: q = 8'h00;
            12'hB38: q = 8'h00;
            12'hB39: q = 8'h00;
            12'hB3A: q = 8'h00;
            12'hB3B: q = 8'h00;
            12'hB3C: q = 8'h00;
            12'hB3D: q = 8'h00;
            12'hB3E: q = 8'h00;
            12'hB3F: q = 8'h00;
            12'hB40: q = 8'h00;
            12'hB41: q = 8'h00;
            12'hB42: q = 8'h00;
            12'hB43: q = 8'h00;
            12'hB44: q = 8'h00;
            12'hB45: q = 8'h00;
            12'hB46: q = 8'h00;
            12'hB47: q = 8'h00;
            12'hB48: q = 8'h00;
            12'hB49: q = 8'h00;
            12'hB4A: q = 8'h00;
            12'hB4B: q = 8'h00;
            12'hB4C: q = 8'h00;
            12'hB4D: q = 8'h00;
            12'hB4E: q = 8'h00;
            12'hB4F: q = 8'h00;
            12'hB50: q = 8'h00;
            12'hB51: q = 8'h00;
            12'hB52: q = 8'h00;
            12'hB53: q = 8'h00;
            12'hB54: q = 8'h00;
            12'hB55: q = 8'h00;
            12'hB56: q = 8'h00;
            12'hB57: q = 8'h00;
            12'hB58: q = 8'h00;
            12'hB59: q = 8'h00;
            12'hB5A: q = 8'h00;
            12'hB5B: q = 8'h00;
            12'hB5C: q = 8'h00;
            12'hB5D: q = 8'h00;
            12'hB5E: q = 8'h00;
            12'hB5F: q = 8'h00;
            12'hB60: q = 8'h00;
            12'hB61: q = 8'h00;
            12'hB62: q = 8'h00;
            12'hB63: q = 8'h00;
            12'hB64: q = 8'h00;
            12'hB65: q = 8'h00;
            12'hB66: q = 8'h00;
            12'hB67: q = 8'h00;
            12'hB68: q = 8'h00;
            12'hB69: q = 8'h00;
            12'hB6A: q = 8'h00;
            12'hB6B: q = 8'h00;
            12'hB6C: q = 8'h00;
            12'hB6D: q = 8'h00;
            12'hB6E: q = 8'h00;
            12'hB6F: q = 8'h00;
            12'hB70: q = 8'h00;
            12'hB71: q = 8'h00;
            12'hB72: q = 8'h00;
            12'hB73: q = 8'h00;
            12'hB74: q = 8'h00;
            12'hB75: q = 8'h00;
            12'hB76: q = 8'h00;
            12'hB77: q = 8'h00;
            12'hB78: q = 8'h00;
            12'hB79: q = 8'h00;
            12'hB7A: q = 8'h00;
            12'hB7B: q = 8'h00;
            12'hB7C: q = 8'h00;
            12'hB7D: q = 8'h00;
            12'hB7E: q = 8'h00;
            12'hB7F: q = 8'h00;
            12'hB80: q = 8'h00;
            12'hB81: q = 8'h00;
            12'hB82: q = 8'h00;
            12'hB83: q = 8'h00;
            12'hB84: q = 8'h00;
            12'hB85: q = 8'h00;
            12'hB86: q = 8'h00;
            12'hB87: q = 8'h00;
            12'hB88: q = 8'h00;
            12'hB89: q = 8'h00;
            12'hB8A: q = 8'h00;
            12'hB8B: q = 8'h00;
            12'hB8C: q = 8'h00;
            12'hB8D: q = 8'h00;
            12'hB8E: q = 8'h00;
            12'hB8F: q = 8'h00;
            12'hB90: q = 8'h00;
            12'hB91: q = 8'h00;
            12'hB92: q = 8'h00;
            12'hB93: q = 8'h00;
            12'hB94: q = 8'h00;
            12'hB95: q = 8'h00;
            12'hB96: q = 8'h00;
            12'hB97: q = 8'h00;
            12'hB98: q = 8'h00;
            12'hB99: q = 8'h00;
            12'hB9A: q = 8'h00;
            12'hB9B: q = 8'h00;
            12'hB9C: q = 8'h00;
            12'hB9D: q = 8'h00;
            12'hB9E: q = 8'h00;
            12'hB9F: q = 8'h00;
            12'hBA0: q = 8'h00;
            12'hBA1: q = 8'h00;
            12'hBA2: q = 8'h00;
            12'hBA3: q = 8'h00;
            12'hBA4: q = 8'h00;
            12'hBA5: q = 8'h00;
            12'hBA6: q = 8'h00;
            12'hBA7: q = 8'h00;
            12'hBA8: q = 8'h00;
            12'hBA9: q = 8'h00;
            12'hBAA: q = 8'h00;
            12'hBAB: q = 8'h00;
            12'hBAC: q = 8'h00;
            12'hBAD: q = 8'h00;
            12'hBAE: q = 8'h00;
            12'hBAF: q = 8'h00;
            12'hBB0: q = 8'h00;
            12'hBB1: q = 8'h00;
            12'hBB2: q = 8'h00;
            12'hBB3: q = 8'h00;
            12'hBB4: q = 8'h00;
            12'hBB5: q = 8'h00;
            12'hBB6: q = 8'h00;
            12'hBB7: q = 8'h00;
            12'hBB8: q = 8'h00;
            12'hBB9: q = 8'h00;
            12'hBBA: q = 8'h00;
            12'hBBB: q = 8'h00;
            12'hBBC: q = 8'h00;
            12'hBBD: q = 8'h00;
            12'hBBE: q = 8'h00;
            12'hBBF: q = 8'h00;
            12'hBC0: q = 8'h00;
            12'hBC1: q = 8'h00;
            12'hBC2: q = 8'h00;
            12'hBC3: q = 8'h00;
            12'hBC4: q = 8'h00;
            12'hBC5: q = 8'h00;
            12'hBC6: q = 8'h00;
            12'hBC7: q = 8'h00;
            12'hBC8: q = 8'h00;
            12'hBC9: q = 8'h00;
            12'hBCA: q = 8'h00;
            12'hBCB: q = 8'h00;
            12'hBCC: q = 8'h00;
            12'hBCD: q = 8'h00;
            12'hBCE: q = 8'h00;
            12'hBCF: q = 8'h00;
            12'hBD0: q = 8'h00;
            12'hBD1: q = 8'h00;
            12'hBD2: q = 8'h00;
            12'hBD3: q = 8'h00;
            12'hBD4: q = 8'h00;
            12'hBD5: q = 8'h00;
            12'hBD6: q = 8'h00;
            12'hBD7: q = 8'h00;
            12'hBD8: q = 8'h00;
            12'hBD9: q = 8'h00;
            12'hBDA: q = 8'h00;
            12'hBDB: q = 8'h00;
            12'hBDC: q = 8'h00;
            12'hBDD: q = 8'h00;
            12'hBDE: q = 8'h00;
            12'hBDF: q = 8'h00;
            12'hBE0: q = 8'h00;
            12'hBE1: q = 8'h00;
            12'hBE2: q = 8'h00;
            12'hBE3: q = 8'h00;
            12'hBE4: q = 8'h00;
            12'hBE5: q = 8'h00;
            12'hBE6: q = 8'h00;
            12'hBE7: q = 8'h00;
            12'hBE8: q = 8'h00;
            12'hBE9: q = 8'h00;
            12'hBEA: q = 8'h00;
            12'hBEB: q = 8'h00;
            12'hBEC: q = 8'h00;
            12'hBED: q = 8'h00;
            12'hBEE: q = 8'h00;
            12'hBEF: q = 8'h00;
            12'hBF0: q = 8'h00;
            12'hBF1: q = 8'h00;
            12'hBF2: q = 8'h00;
            12'hBF3: q = 8'h00;
            12'hBF4: q = 8'h00;
            12'hBF5: q = 8'h00;
            12'hBF6: q = 8'h00;
            12'hBF7: q = 8'h00;
            12'hBF8: q = 8'h00;
            12'hBF9: q = 8'h00;
            12'hBFA: q = 8'h00;
            12'hBFB: q = 8'h00;
            12'hBFC: q = 8'h00;
            12'hBFD: q = 8'h00;
            12'hBFE: q = 8'h00;
            12'hBFF: q = 8'h00;
            12'hC00: q = 8'h00;
            12'hC01: q = 8'h00;
            12'hC02: q = 8'h00;
            12'hC03: q = 8'h00;
            12'hC04: q = 8'h00;
            12'hC05: q = 8'h00;
            12'hC06: q = 8'h00;
            12'hC07: q = 8'h00;
            12'hC08: q = 8'h00;
            12'hC09: q = 8'h00;
            12'hC0A: q = 8'h00;
            12'hC0B: q = 8'h00;
            12'hC0C: q = 8'h00;
            12'hC0D: q = 8'h00;
            12'hC0E: q = 8'h00;
            12'hC0F: q = 8'h00;
            12'hC10: q = 8'h00;
            12'hC11: q = 8'h00;
            12'hC12: q = 8'h00;
            12'hC13: q = 8'h00;
            12'hC14: q = 8'h00;
            12'hC15: q = 8'h00;
            12'hC16: q = 8'h00;
            12'hC17: q = 8'h00;
            12'hC18: q = 8'h00;
            12'hC19: q = 8'h00;
            12'hC1A: q = 8'h00;
            12'hC1B: q = 8'h00;
            12'hC1C: q = 8'h00;
            12'hC1D: q = 8'h00;
            12'hC1E: q = 8'h00;
            12'hC1F: q = 8'h00;
            12'hC20: q = 8'h00;
            12'hC21: q = 8'h00;
            12'hC22: q = 8'h00;
            12'hC23: q = 8'h00;
            12'hC24: q = 8'h00;
            12'hC25: q = 8'h00;
            12'hC26: q = 8'h00;
            12'hC27: q = 8'h00;
            12'hC28: q = 8'h00;
            12'hC29: q = 8'h00;
            12'hC2A: q = 8'h00;
            12'hC2B: q = 8'h00;
            12'hC2C: q = 8'h00;
            12'hC2D: q = 8'h00;
            12'hC2E: q = 8'h00;
            12'hC2F: q = 8'h00;
            12'hC30: q = 8'h00;
            12'hC31: q = 8'h00;
            12'hC32: q = 8'h00;
            12'hC33: q = 8'h00;
            12'hC34: q = 8'h00;
            12'hC35: q = 8'h00;
            12'hC36: q = 8'h00;
            12'hC37: q = 8'h00;
            12'hC38: q = 8'h00;
            12'hC39: q = 8'h00;
            12'hC3A: q = 8'h00;
            12'hC3B: q = 8'h00;
            12'hC3C: q = 8'h00;
            12'hC3D: q = 8'h00;
            12'hC3E: q = 8'h00;
            12'hC3F: q = 8'h00;
            12'hC40: q = 8'h00;
            12'hC41: q = 8'h00;
            12'hC42: q = 8'h00;
            12'hC43: q = 8'h00;
            12'hC44: q = 8'h00;
            12'hC45: q = 8'h00;
            12'hC46: q = 8'h00;
            12'hC47: q = 8'h00;
            12'hC48: q = 8'h00;
            12'hC49: q = 8'h00;
            12'hC4A: q = 8'h00;
            12'hC4B: q = 8'h00;
            12'hC4C: q = 8'h00;
            12'hC4D: q = 8'h00;
            12'hC4E: q = 8'h00;
            12'hC4F: q = 8'h00;
            12'hC50: q = 8'h00;
            12'hC51: q = 8'h00;
            12'hC52: q = 8'h00;
            12'hC53: q = 8'h00;
            12'hC54: q = 8'h00;
            12'hC55: q = 8'h00;
            12'hC56: q = 8'h00;
            12'hC57: q = 8'h00;
            12'hC58: q = 8'h00;
            12'hC59: q = 8'h00;
            12'hC5A: q = 8'h00;
            12'hC5B: q = 8'h00;
            12'hC5C: q = 8'h00;
            12'hC5D: q = 8'h00;
            12'hC5E: q = 8'h00;
            12'hC5F: q = 8'h00;
            12'hC60: q = 8'h00;
            12'hC61: q = 8'h00;
            12'hC62: q = 8'h00;
            12'hC63: q = 8'h00;
            12'hC64: q = 8'h00;
            12'hC65: q = 8'h00;
            12'hC66: q = 8'h00;
            12'hC67: q = 8'h00;
            12'hC68: q = 8'h00;
            12'hC69: q = 8'h00;
            12'hC6A: q = 8'h00;
            12'hC6B: q = 8'h00;
            12'hC6C: q = 8'h00;
            12'hC6D: q = 8'h00;
            12'hC6E: q = 8'h00;
            12'hC6F: q = 8'h00;
            12'hC70: q = 8'h00;
            12'hC71: q = 8'h00;
            12'hC72: q = 8'h00;
            12'hC73: q = 8'h00;
            12'hC74: q = 8'h00;
            12'hC75: q = 8'h00;
            12'hC76: q = 8'h00;
            12'hC77: q = 8'h00;
            12'hC78: q = 8'h00;
            12'hC79: q = 8'h00;
            12'hC7A: q = 8'h00;
            12'hC7B: q = 8'h00;
            12'hC7C: q = 8'h00;
            12'hC7D: q = 8'h00;
            12'hC7E: q = 8'h00;
            12'hC7F: q = 8'h00;
            12'hC80: q = 8'h00;
            12'hC81: q = 8'h00;
            12'hC82: q = 8'h00;
            12'hC83: q = 8'h00;
            12'hC84: q = 8'h00;
            12'hC85: q = 8'h00;
            12'hC86: q = 8'h00;
            12'hC87: q = 8'h00;
            12'hC88: q = 8'h00;
            12'hC89: q = 8'h00;
            12'hC8A: q = 8'h00;
            12'hC8B: q = 8'h00;
            12'hC8C: q = 8'h00;
            12'hC8D: q = 8'h00;
            12'hC8E: q = 8'h00;
            12'hC8F: q = 8'h00;
            12'hC90: q = 8'h00;
            12'hC91: q = 8'h00;
            12'hC92: q = 8'h00;
            12'hC93: q = 8'h00;
            12'hC94: q = 8'h00;
            12'hC95: q = 8'h00;
            12'hC96: q = 8'h00;
            12'hC97: q = 8'h00;
            12'hC98: q = 8'h00;
            12'hC99: q = 8'h00;
            12'hC9A: q = 8'h00;
            12'hC9B: q = 8'h00;
            12'hC9C: q = 8'h00;
            12'hC9D: q = 8'h00;
            12'hC9E: q = 8'h00;
            12'hC9F: q = 8'h00;
            12'hCA0: q = 8'h00;
            12'hCA1: q = 8'h00;
            12'hCA2: q = 8'h00;
            12'hCA3: q = 8'h00;
            12'hCA4: q = 8'h00;
            12'hCA5: q = 8'h00;
            12'hCA6: q = 8'h00;
            12'hCA7: q = 8'h00;
            12'hCA8: q = 8'h00;
            12'hCA9: q = 8'h00;
            12'hCAA: q = 8'h00;
            12'hCAB: q = 8'h00;
            12'hCAC: q = 8'h00;
            12'hCAD: q = 8'h00;
            12'hCAE: q = 8'h00;
            12'hCAF: q = 8'h00;
            12'hCB0: q = 8'h00;
            12'hCB1: q = 8'h00;
            12'hCB2: q = 8'h00;
            12'hCB3: q = 8'h00;
            12'hCB4: q = 8'h00;
            12'hCB5: q = 8'h00;
            12'hCB6: q = 8'h00;
            12'hCB7: q = 8'h00;
            12'hCB8: q = 8'h00;
            12'hCB9: q = 8'h00;
            12'hCBA: q = 8'h00;
            12'hCBB: q = 8'h00;
            12'hCBC: q = 8'h00;
            12'hCBD: q = 8'h00;
            12'hCBE: q = 8'h00;
            12'hCBF: q = 8'h00;
            12'hCC0: q = 8'h00;
            12'hCC1: q = 8'h00;
            12'hCC2: q = 8'h00;
            12'hCC3: q = 8'h00;
            12'hCC4: q = 8'h00;
            12'hCC5: q = 8'h00;
            12'hCC6: q = 8'h00;
            12'hCC7: q = 8'h00;
            12'hCC8: q = 8'h00;
            12'hCC9: q = 8'h00;
            12'hCCA: q = 8'h00;
            12'hCCB: q = 8'h00;
            12'hCCC: q = 8'h00;
            12'hCCD: q = 8'h00;
            12'hCCE: q = 8'h00;
            12'hCCF: q = 8'h00;
            12'hCD0: q = 8'h00;
            12'hCD1: q = 8'h00;
            12'hCD2: q = 8'h00;
            12'hCD3: q = 8'h00;
            12'hCD4: q = 8'h00;
            12'hCD5: q = 8'h00;
            12'hCD6: q = 8'h00;
            12'hCD7: q = 8'h00;
            12'hCD8: q = 8'h00;
            12'hCD9: q = 8'h00;
            12'hCDA: q = 8'h00;
            12'hCDB: q = 8'h00;
            12'hCDC: q = 8'h00;
            12'hCDD: q = 8'h00;
            12'hCDE: q = 8'h00;
            12'hCDF: q = 8'h00;
            12'hCE0: q = 8'h00;
            12'hCE1: q = 8'h00;
            12'hCE2: q = 8'h00;
            12'hCE3: q = 8'h00;
            12'hCE4: q = 8'h00;
            12'hCE5: q = 8'h00;
            12'hCE6: q = 8'h00;
            12'hCE7: q = 8'h00;
            12'hCE8: q = 8'h00;
            12'hCE9: q = 8'h00;
            12'hCEA: q = 8'h00;
            12'hCEB: q = 8'h00;
            12'hCEC: q = 8'h00;
            12'hCED: q = 8'h00;
            12'hCEE: q = 8'h00;
            12'hCEF: q = 8'h00;
            12'hCF0: q = 8'h00;
            12'hCF1: q = 8'h00;
            12'hCF2: q = 8'h00;
            12'hCF3: q = 8'h00;
            12'hCF4: q = 8'h00;
            12'hCF5: q = 8'h00;
            12'hCF6: q = 8'h00;
            12'hCF7: q = 8'h00;
            12'hCF8: q = 8'h00;
            12'hCF9: q = 8'h00;
            12'hCFA: q = 8'h00;
            12'hCFB: q = 8'h00;
            12'hCFC: q = 8'h00;
            12'hCFD: q = 8'h00;
            12'hCFE: q = 8'h00;
            12'hCFF: q = 8'h00;
            12'hD00: q = 8'h00;
            12'hD01: q = 8'h00;
            12'hD02: q = 8'h00;
            12'hD03: q = 8'h00;
            12'hD04: q = 8'h00;
            12'hD05: q = 8'h00;
            12'hD06: q = 8'h00;
            12'hD07: q = 8'h00;
            12'hD08: q = 8'h00;
            12'hD09: q = 8'h00;
            12'hD0A: q = 8'h00;
            12'hD0B: q = 8'h00;
            12'hD0C: q = 8'h00;
            12'hD0D: q = 8'h00;
            12'hD0E: q = 8'h00;
            12'hD0F: q = 8'h00;
            12'hD10: q = 8'h00;
            12'hD11: q = 8'h00;
            12'hD12: q = 8'h00;
            12'hD13: q = 8'h00;
            12'hD14: q = 8'h00;
            12'hD15: q = 8'h00;
            12'hD16: q = 8'h00;
            12'hD17: q = 8'h00;
            12'hD18: q = 8'h00;
            12'hD19: q = 8'h00;
            12'hD1A: q = 8'h00;
            12'hD1B: q = 8'h00;
            12'hD1C: q = 8'h00;
            12'hD1D: q = 8'h00;
            12'hD1E: q = 8'h00;
            12'hD1F: q = 8'h00;
            12'hD20: q = 8'h00;
            12'hD21: q = 8'h00;
            12'hD22: q = 8'h00;
            12'hD23: q = 8'h00;
            12'hD24: q = 8'h00;
            12'hD25: q = 8'h00;
            12'hD26: q = 8'h00;
            12'hD27: q = 8'h00;
            12'hD28: q = 8'h00;
            12'hD29: q = 8'h00;
            12'hD2A: q = 8'h00;
            12'hD2B: q = 8'h00;
            12'hD2C: q = 8'h00;
            12'hD2D: q = 8'h00;
            12'hD2E: q = 8'h00;
            12'hD2F: q = 8'h00;
            12'hD30: q = 8'h00;
            12'hD31: q = 8'h00;
            12'hD32: q = 8'h00;
            12'hD33: q = 8'h00;
            12'hD34: q = 8'h00;
            12'hD35: q = 8'h00;
            12'hD36: q = 8'h00;
            12'hD37: q = 8'h00;
            12'hD38: q = 8'h00;
            12'hD39: q = 8'h00;
            12'hD3A: q = 8'h00;
            12'hD3B: q = 8'h00;
            12'hD3C: q = 8'h00;
            12'hD3D: q = 8'h00;
            12'hD3E: q = 8'h00;
            12'hD3F: q = 8'h00;
            12'hD40: q = 8'h00;
            12'hD41: q = 8'h00;
            12'hD42: q = 8'h00;
            12'hD43: q = 8'h00;
            12'hD44: q = 8'h00;
            12'hD45: q = 8'h00;
            12'hD46: q = 8'h00;
            12'hD47: q = 8'h00;
            12'hD48: q = 8'h00;
            12'hD49: q = 8'h00;
            12'hD4A: q = 8'h00;
            12'hD4B: q = 8'h00;
            12'hD4C: q = 8'h00;
            12'hD4D: q = 8'h00;
            12'hD4E: q = 8'h00;
            12'hD4F: q = 8'h00;
            12'hD50: q = 8'h00;
            12'hD51: q = 8'h00;
            12'hD52: q = 8'h00;
            12'hD53: q = 8'h00;
            12'hD54: q = 8'h00;
            12'hD55: q = 8'h00;
            12'hD56: q = 8'h00;
            12'hD57: q = 8'h00;
            12'hD58: q = 8'h00;
            12'hD59: q = 8'h00;
            12'hD5A: q = 8'h00;
            12'hD5B: q = 8'h00;
            12'hD5C: q = 8'h00;
            12'hD5D: q = 8'h00;
            12'hD5E: q = 8'h00;
            12'hD5F: q = 8'h00;
            12'hD60: q = 8'h00;
            12'hD61: q = 8'h00;
            12'hD62: q = 8'h00;
            12'hD63: q = 8'h00;
            12'hD64: q = 8'h00;
            12'hD65: q = 8'h00;
            12'hD66: q = 8'h00;
            12'hD67: q = 8'h00;
            12'hD68: q = 8'h00;
            12'hD69: q = 8'h00;
            12'hD6A: q = 8'h00;
            12'hD6B: q = 8'h00;
            12'hD6C: q = 8'h00;
            12'hD6D: q = 8'h00;
            12'hD6E: q = 8'h00;
            12'hD6F: q = 8'h00;
            12'hD70: q = 8'h00;
            12'hD71: q = 8'h00;
            12'hD72: q = 8'h00;
            12'hD73: q = 8'h00;
            12'hD74: q = 8'h00;
            12'hD75: q = 8'h00;
            12'hD76: q = 8'h00;
            12'hD77: q = 8'h00;
            12'hD78: q = 8'h00;
            12'hD79: q = 8'h00;
            12'hD7A: q = 8'h00;
            12'hD7B: q = 8'h00;
            12'hD7C: q = 8'h00;
            12'hD7D: q = 8'h00;
            12'hD7E: q = 8'h00;
            12'hD7F: q = 8'h00;
            12'hD80: q = 8'h00;
            12'hD81: q = 8'h00;
            12'hD82: q = 8'h00;
            12'hD83: q = 8'h00;
            12'hD84: q = 8'h00;
            12'hD85: q = 8'h00;
            12'hD86: q = 8'h00;
            12'hD87: q = 8'h00;
            12'hD88: q = 8'h00;
            12'hD89: q = 8'h00;
            12'hD8A: q = 8'h00;
            12'hD8B: q = 8'h00;
            12'hD8C: q = 8'h00;
            12'hD8D: q = 8'h00;
            12'hD8E: q = 8'h00;
            12'hD8F: q = 8'h00;
            12'hD90: q = 8'h00;
            12'hD91: q = 8'h00;
            12'hD92: q = 8'h00;
            12'hD93: q = 8'h00;
            12'hD94: q = 8'h00;
            12'hD95: q = 8'h00;
            12'hD96: q = 8'h00;
            12'hD97: q = 8'h00;
            12'hD98: q = 8'h00;
            12'hD99: q = 8'h00;
            12'hD9A: q = 8'h00;
            12'hD9B: q = 8'h00;
            12'hD9C: q = 8'h00;
            12'hD9D: q = 8'h00;
            12'hD9E: q = 8'h00;
            12'hD9F: q = 8'h00;
            12'hDA0: q = 8'h00;
            12'hDA1: q = 8'h00;
            12'hDA2: q = 8'h00;
            12'hDA3: q = 8'h00;
            12'hDA4: q = 8'h00;
            12'hDA5: q = 8'h00;
            12'hDA6: q = 8'h00;
            12'hDA7: q = 8'h00;
            12'hDA8: q = 8'h00;
            12'hDA9: q = 8'h00;
            12'hDAA: q = 8'h00;
            12'hDAB: q = 8'h00;
            12'hDAC: q = 8'h00;
            12'hDAD: q = 8'h00;
            12'hDAE: q = 8'h00;
            12'hDAF: q = 8'h00;
            12'hDB0: q = 8'h00;
            12'hDB1: q = 8'h00;
            12'hDB2: q = 8'h00;
            12'hDB3: q = 8'h00;
            12'hDB4: q = 8'h00;
            12'hDB5: q = 8'h00;
            12'hDB6: q = 8'h00;
            12'hDB7: q = 8'h00;
            12'hDB8: q = 8'h00;
            12'hDB9: q = 8'h00;
            12'hDBA: q = 8'h00;
            12'hDBB: q = 8'h00;
            12'hDBC: q = 8'h00;
            12'hDBD: q = 8'h00;
            12'hDBE: q = 8'h00;
            12'hDBF: q = 8'h00;
            12'hDC0: q = 8'h00;
            12'hDC1: q = 8'h00;
            12'hDC2: q = 8'h00;
            12'hDC3: q = 8'h00;
            12'hDC4: q = 8'h00;
            12'hDC5: q = 8'h00;
            12'hDC6: q = 8'h00;
            12'hDC7: q = 8'h00;
            12'hDC8: q = 8'h00;
            12'hDC9: q = 8'h00;
            12'hDCA: q = 8'h00;
            12'hDCB: q = 8'h00;
            12'hDCC: q = 8'h00;
            12'hDCD: q = 8'h00;
            12'hDCE: q = 8'h00;
            12'hDCF: q = 8'h00;
            12'hDD0: q = 8'h00;
            12'hDD1: q = 8'h00;
            12'hDD2: q = 8'h00;
            12'hDD3: q = 8'h00;
            12'hDD4: q = 8'h00;
            12'hDD5: q = 8'h00;
            12'hDD6: q = 8'h00;
            12'hDD7: q = 8'h00;
            12'hDD8: q = 8'h00;
            12'hDD9: q = 8'h00;
            12'hDDA: q = 8'h00;
            12'hDDB: q = 8'h00;
            12'hDDC: q = 8'h00;
            12'hDDD: q = 8'h00;
            12'hDDE: q = 8'h00;
            12'hDDF: q = 8'h00;
            12'hDE0: q = 8'h00;
            12'hDE1: q = 8'h00;
            12'hDE2: q = 8'h00;
            12'hDE3: q = 8'h00;
            12'hDE4: q = 8'h00;
            12'hDE5: q = 8'h00;
            12'hDE6: q = 8'h00;
            12'hDE7: q = 8'h00;
            12'hDE8: q = 8'h00;
            12'hDE9: q = 8'h00;
            12'hDEA: q = 8'h00;
            12'hDEB: q = 8'h00;
            12'hDEC: q = 8'h00;
            12'hDED: q = 8'h00;
            12'hDEE: q = 8'h00;
            12'hDEF: q = 8'h00;
            12'hDF0: q = 8'h00;
            12'hDF1: q = 8'h00;
            12'hDF2: q = 8'h00;
            12'hDF3: q = 8'h00;
            12'hDF4: q = 8'h00;
            12'hDF5: q = 8'h00;
            12'hDF6: q = 8'h00;
            12'hDF7: q = 8'h00;
            12'hDF8: q = 8'h00;
            12'hDF9: q = 8'h00;
            12'hDFA: q = 8'h00;
            12'hDFB: q = 8'h00;
            12'hDFC: q = 8'h00;
            12'hDFD: q = 8'h00;
            12'hDFE: q = 8'h00;
            12'hDFF: q = 8'h00;
            12'hE00: q = 8'h00;
            12'hE01: q = 8'h00;
            12'hE02: q = 8'h00;
            12'hE03: q = 8'h00;
            12'hE04: q = 8'h00;
            12'hE05: q = 8'h00;
            12'hE06: q = 8'h00;
            12'hE07: q = 8'h00;
            12'hE08: q = 8'h00;
            12'hE09: q = 8'h00;
            12'hE0A: q = 8'h00;
            12'hE0B: q = 8'h00;
            12'hE0C: q = 8'h00;
            12'hE0D: q = 8'h00;
            12'hE0E: q = 8'h00;
            12'hE0F: q = 8'h00;
            12'hE10: q = 8'h00;
            12'hE11: q = 8'h00;
            12'hE12: q = 8'h00;
            12'hE13: q = 8'h00;
            12'hE14: q = 8'h00;
            12'hE15: q = 8'h00;
            12'hE16: q = 8'h00;
            12'hE17: q = 8'h00;
            12'hE18: q = 8'h00;
            12'hE19: q = 8'h00;
            12'hE1A: q = 8'h00;
            12'hE1B: q = 8'h00;
            12'hE1C: q = 8'h00;
            12'hE1D: q = 8'h00;
            12'hE1E: q = 8'h00;
            12'hE1F: q = 8'h00;
            12'hE20: q = 8'h00;
            12'hE21: q = 8'h00;
            12'hE22: q = 8'h00;
            12'hE23: q = 8'h00;
            12'hE24: q = 8'h00;
            12'hE25: q = 8'h00;
            12'hE26: q = 8'h00;
            12'hE27: q = 8'h00;
            12'hE28: q = 8'h00;
            12'hE29: q = 8'h00;
            12'hE2A: q = 8'h00;
            12'hE2B: q = 8'h00;
            12'hE2C: q = 8'h00;
            12'hE2D: q = 8'h00;
            12'hE2E: q = 8'h00;
            12'hE2F: q = 8'h00;
            12'hE30: q = 8'h00;
            12'hE31: q = 8'h00;
            12'hE32: q = 8'h00;
            12'hE33: q = 8'h00;
            12'hE34: q = 8'h00;
            12'hE35: q = 8'h00;
            12'hE36: q = 8'h00;
            12'hE37: q = 8'h00;
            12'hE38: q = 8'h00;
            12'hE39: q = 8'h00;
            12'hE3A: q = 8'h00;
            12'hE3B: q = 8'h00;
            12'hE3C: q = 8'h00;
            12'hE3D: q = 8'h00;
            12'hE3E: q = 8'h00;
            12'hE3F: q = 8'h00;
            12'hE40: q = 8'h00;
            12'hE41: q = 8'h00;
            12'hE42: q = 8'h00;
            12'hE43: q = 8'h00;
            12'hE44: q = 8'h00;
            12'hE45: q = 8'h00;
            12'hE46: q = 8'h00;
            12'hE47: q = 8'h00;
            12'hE48: q = 8'h00;
            12'hE49: q = 8'h00;
            12'hE4A: q = 8'h00;
            12'hE4B: q = 8'h00;
            12'hE4C: q = 8'h00;
            12'hE4D: q = 8'h00;
            12'hE4E: q = 8'h00;
            12'hE4F: q = 8'h00;
            12'hE50: q = 8'h00;
            12'hE51: q = 8'h00;
            12'hE52: q = 8'h00;
            12'hE53: q = 8'h00;
            12'hE54: q = 8'h00;
            12'hE55: q = 8'h00;
            12'hE56: q = 8'h00;
            12'hE57: q = 8'h00;
            12'hE58: q = 8'h00;
            12'hE59: q = 8'h00;
            12'hE5A: q = 8'h00;
            12'hE5B: q = 8'h00;
            12'hE5C: q = 8'h00;
            12'hE5D: q = 8'h00;
            12'hE5E: q = 8'h00;
            12'hE5F: q = 8'h00;
            12'hE60: q = 8'h00;
            12'hE61: q = 8'h00;
            12'hE62: q = 8'h00;
            12'hE63: q = 8'h00;
            12'hE64: q = 8'h00;
            12'hE65: q = 8'h00;
            12'hE66: q = 8'h00;
            12'hE67: q = 8'h00;
            12'hE68: q = 8'h00;
            12'hE69: q = 8'h00;
            12'hE6A: q = 8'h00;
            12'hE6B: q = 8'h00;
            12'hE6C: q = 8'h00;
            12'hE6D: q = 8'h00;
            12'hE6E: q = 8'h00;
            12'hE6F: q = 8'h00;
            12'hE70: q = 8'h00;
            12'hE71: q = 8'h00;
            12'hE72: q = 8'h00;
            12'hE73: q = 8'h00;
            12'hE74: q = 8'h00;
            12'hE75: q = 8'h00;
            12'hE76: q = 8'h00;
            12'hE77: q = 8'h00;
            12'hE78: q = 8'h00;
            12'hE79: q = 8'h00;
            12'hE7A: q = 8'h00;
            12'hE7B: q = 8'h00;
            12'hE7C: q = 8'h00;
            12'hE7D: q = 8'h00;
            12'hE7E: q = 8'h00;
            12'hE7F: q = 8'h00;
            12'hE80: q = 8'h00;
            12'hE81: q = 8'h00;
            12'hE82: q = 8'h00;
            12'hE83: q = 8'h00;
            12'hE84: q = 8'h00;
            12'hE85: q = 8'h00;
            12'hE86: q = 8'h00;
            12'hE87: q = 8'h00;
            12'hE88: q = 8'h00;
            12'hE89: q = 8'h00;
            12'hE8A: q = 8'h00;
            12'hE8B: q = 8'h00;
            12'hE8C: q = 8'h00;
            12'hE8D: q = 8'h00;
            12'hE8E: q = 8'h00;
            12'hE8F: q = 8'h00;
            12'hE90: q = 8'h00;
            12'hE91: q = 8'h00;
            12'hE92: q = 8'h00;
            12'hE93: q = 8'h00;
            12'hE94: q = 8'h00;
            12'hE95: q = 8'h00;
            12'hE96: q = 8'h00;
            12'hE97: q = 8'h00;
            12'hE98: q = 8'h00;
            12'hE99: q = 8'h00;
            12'hE9A: q = 8'h00;
            12'hE9B: q = 8'h00;
            12'hE9C: q = 8'h00;
            12'hE9D: q = 8'h00;
            12'hE9E: q = 8'h00;
            12'hE9F: q = 8'h00;
            12'hEA0: q = 8'h00;
            12'hEA1: q = 8'h00;
            12'hEA2: q = 8'h00;
            12'hEA3: q = 8'h00;
            12'hEA4: q = 8'h00;
            12'hEA5: q = 8'h00;
            12'hEA6: q = 8'h00;
            12'hEA7: q = 8'h00;
            12'hEA8: q = 8'h00;
            12'hEA9: q = 8'h00;
            12'hEAA: q = 8'h00;
            12'hEAB: q = 8'h00;
            12'hEAC: q = 8'h00;
            12'hEAD: q = 8'h00;
            12'hEAE: q = 8'h00;
            12'hEAF: q = 8'h00;
            12'hEB0: q = 8'h00;
            12'hEB1: q = 8'h00;
            12'hEB2: q = 8'h00;
            12'hEB3: q = 8'h00;
            12'hEB4: q = 8'h00;
            12'hEB5: q = 8'h00;
            12'hEB6: q = 8'h00;
            12'hEB7: q = 8'h00;
            12'hEB8: q = 8'h00;
            12'hEB9: q = 8'h00;
            12'hEBA: q = 8'h00;
            12'hEBB: q = 8'h00;
            12'hEBC: q = 8'h00;
            12'hEBD: q = 8'h00;
            12'hEBE: q = 8'h00;
            12'hEBF: q = 8'h00;
            12'hEC0: q = 8'h00;
            12'hEC1: q = 8'h00;
            12'hEC2: q = 8'h00;
            12'hEC3: q = 8'h00;
            12'hEC4: q = 8'h00;
            12'hEC5: q = 8'h00;
            12'hEC6: q = 8'h00;
            12'hEC7: q = 8'h00;
            12'hEC8: q = 8'h00;
            12'hEC9: q = 8'h00;
            12'hECA: q = 8'h00;
            12'hECB: q = 8'h00;
            12'hECC: q = 8'h00;
            12'hECD: q = 8'h00;
            12'hECE: q = 8'h00;
            12'hECF: q = 8'h00;
            12'hED0: q = 8'h00;
            12'hED1: q = 8'h00;
            12'hED2: q = 8'h00;
            12'hED3: q = 8'h00;
            12'hED4: q = 8'h00;
            12'hED5: q = 8'h00;
            12'hED6: q = 8'h00;
            12'hED7: q = 8'h00;
            12'hED8: q = 8'h00;
            12'hED9: q = 8'h00;
            12'hEDA: q = 8'h00;
            12'hEDB: q = 8'h00;
            12'hEDC: q = 8'h00;
            12'hEDD: q = 8'h00;
            12'hEDE: q = 8'h00;
            12'hEDF: q = 8'h00;
            12'hEE0: q = 8'h00;
            12'hEE1: q = 8'h00;
            12'hEE2: q = 8'h00;
            12'hEE3: q = 8'h00;
            12'hEE4: q = 8'h00;
            12'hEE5: q = 8'h00;
            12'hEE6: q = 8'h00;
            12'hEE7: q = 8'h00;
            12'hEE8: q = 8'h00;
            12'hEE9: q = 8'h00;
            12'hEEA: q = 8'h00;
            12'hEEB: q = 8'h00;
            12'hEEC: q = 8'h00;
            12'hEED: q = 8'h00;
            12'hEEE: q = 8'h00;
            12'hEEF: q = 8'h00;
            12'hEF0: q = 8'h00;
            12'hEF1: q = 8'h00;
            12'hEF2: q = 8'h00;
            12'hEF3: q = 8'h00;
            12'hEF4: q = 8'h00;
            12'hEF5: q = 8'h00;
            12'hEF6: q = 8'h00;
            12'hEF7: q = 8'h00;
            12'hEF8: q = 8'h00;
            12'hEF9: q = 8'h00;
            12'hEFA: q = 8'h00;
            12'hEFB: q = 8'h00;
            12'hEFC: q = 8'h00;
            12'hEFD: q = 8'h00;
            12'hEFE: q = 8'h00;
            12'hEFF: q = 8'h00;
            12'hF00: q = 8'h00;
            12'hF01: q = 8'h00;
            12'hF02: q = 8'h00;
            12'hF03: q = 8'h00;
            12'hF04: q = 8'h00;
            12'hF05: q = 8'h00;
            12'hF06: q = 8'h00;
            12'hF07: q = 8'h00;
            12'hF08: q = 8'h00;
            12'hF09: q = 8'h00;
            12'hF0A: q = 8'h00;
            12'hF0B: q = 8'h00;
            12'hF0C: q = 8'h00;
            12'hF0D: q = 8'h00;
            12'hF0E: q = 8'h00;
            12'hF0F: q = 8'h00;
            12'hF10: q = 8'h00;
            12'hF11: q = 8'h00;
            12'hF12: q = 8'h00;
            12'hF13: q = 8'h00;
            12'hF14: q = 8'h00;
            12'hF15: q = 8'h00;
            12'hF16: q = 8'h00;
            12'hF17: q = 8'h00;
            12'hF18: q = 8'h00;
            12'hF19: q = 8'h00;
            12'hF1A: q = 8'h00;
            12'hF1B: q = 8'h00;
            12'hF1C: q = 8'h00;
            12'hF1D: q = 8'h00;
            12'hF1E: q = 8'h00;
            12'hF1F: q = 8'h00;
            12'hF20: q = 8'h00;
            12'hF21: q = 8'h00;
            12'hF22: q = 8'h00;
            12'hF23: q = 8'h00;
            12'hF24: q = 8'h00;
            12'hF25: q = 8'h00;
            12'hF26: q = 8'h00;
            12'hF27: q = 8'h00;
            12'hF28: q = 8'h00;
            12'hF29: q = 8'h00;
            12'hF2A: q = 8'h00;
            12'hF2B: q = 8'h00;
            12'hF2C: q = 8'h00;
            12'hF2D: q = 8'h00;
            12'hF2E: q = 8'h00;
            12'hF2F: q = 8'h00;
            12'hF30: q = 8'h00;
            12'hF31: q = 8'h00;
            12'hF32: q = 8'h00;
            12'hF33: q = 8'h00;
            12'hF34: q = 8'h00;
            12'hF35: q = 8'h00;
            12'hF36: q = 8'h00;
            12'hF37: q = 8'h00;
            12'hF38: q = 8'h00;
            12'hF39: q = 8'h00;
            12'hF3A: q = 8'h00;
            12'hF3B: q = 8'h00;
            12'hF3C: q = 8'h00;
            12'hF3D: q = 8'h00;
            12'hF3E: q = 8'h00;
            12'hF3F: q = 8'h00;
            12'hF40: q = 8'h00;
            12'hF41: q = 8'h00;
            12'hF42: q = 8'h00;
            12'hF43: q = 8'h00;
            12'hF44: q = 8'h00;
            12'hF45: q = 8'h00;
            12'hF46: q = 8'h00;
            12'hF47: q = 8'h00;
            12'hF48: q = 8'h00;
            12'hF49: q = 8'h00;
            12'hF4A: q = 8'h00;
            12'hF4B: q = 8'h00;
            12'hF4C: q = 8'h00;
            12'hF4D: q = 8'h00;
            12'hF4E: q = 8'h00;
            12'hF4F: q = 8'h00;
            12'hF50: q = 8'h00;
            12'hF51: q = 8'h00;
            12'hF52: q = 8'h00;
            12'hF53: q = 8'h00;
            12'hF54: q = 8'h00;
            12'hF55: q = 8'h00;
            12'hF56: q = 8'h00;
            12'hF57: q = 8'h00;
            12'hF58: q = 8'h00;
            12'hF59: q = 8'h00;
            12'hF5A: q = 8'h00;
            12'hF5B: q = 8'h00;
            12'hF5C: q = 8'h00;
            12'hF5D: q = 8'h00;
            12'hF5E: q = 8'h00;
            12'hF5F: q = 8'h00;
            12'hF60: q = 8'h00;
            12'hF61: q = 8'h00;
            12'hF62: q = 8'h00;
            12'hF63: q = 8'h00;
            12'hF64: q = 8'h00;
            12'hF65: q = 8'h00;
            12'hF66: q = 8'h00;
            12'hF67: q = 8'h00;
            12'hF68: q = 8'h00;
            12'hF69: q = 8'h00;
            12'hF6A: q = 8'h00;
            12'hF6B: q = 8'h00;
            12'hF6C: q = 8'h00;
            12'hF6D: q = 8'h00;
            12'hF6E: q = 8'h00;
            12'hF6F: q = 8'h00;
            12'hF70: q = 8'h00;
            12'hF71: q = 8'h00;
            12'hF72: q = 8'h00;
            12'hF73: q = 8'h00;
            12'hF74: q = 8'h00;
            12'hF75: q = 8'h00;
            12'hF76: q = 8'h00;
            12'hF77: q = 8'h00;
            12'hF78: q = 8'h00;
            12'hF79: q = 8'h00;
            12'hF7A: q = 8'h00;
            12'hF7B: q = 8'h00;
            12'hF7C: q = 8'h00;
            12'hF7D: q = 8'h00;
            12'hF7E: q = 8'h00;
            12'hF7F: q = 8'h00;
            12'hF80: q = 8'h00;
            12'hF81: q = 8'h00;
            12'hF82: q = 8'h00;
            12'hF83: q = 8'h00;
            12'hF84: q = 8'h00;
            12'hF85: q = 8'h00;
            12'hF86: q = 8'h00;
            12'hF87: q = 8'h00;
            12'hF88: q = 8'h00;
            12'hF89: q = 8'h00;
            12'hF8A: q = 8'h00;
            12'hF8B: q = 8'h00;
            12'hF8C: q = 8'h00;
            12'hF8D: q = 8'h00;
            12'hF8E: q = 8'h00;
            12'hF8F: q = 8'h00;
            12'hF90: q = 8'h00;
            12'hF91: q = 8'h00;
            12'hF92: q = 8'h00;
            12'hF93: q = 8'h00;
            12'hF94: q = 8'h00;
            12'hF95: q = 8'h00;
            12'hF96: q = 8'h00;
            12'hF97: q = 8'h00;
            12'hF98: q = 8'h00;
            12'hF99: q = 8'h00;
            12'hF9A: q = 8'h00;
            12'hF9B: q = 8'h00;
            12'hF9C: q = 8'h00;
            12'hF9D: q = 8'h00;
            12'hF9E: q = 8'h00;
            12'hF9F: q = 8'h00;
            12'hFA0: q = 8'h00;
            12'hFA1: q = 8'h00;
            12'hFA2: q = 8'h00;
            12'hFA3: q = 8'h00;
            12'hFA4: q = 8'h00;
            12'hFA5: q = 8'h00;
            12'hFA6: q = 8'h00;
            12'hFA7: q = 8'h00;
            12'hFA8: q = 8'h00;
            12'hFA9: q = 8'h00;
            12'hFAA: q = 8'h00;
            12'hFAB: q = 8'h00;
            12'hFAC: q = 8'h00;
            12'hFAD: q = 8'h00;
            12'hFAE: q = 8'h00;
            12'hFAF: q = 8'h00;
            12'hFB0: q = 8'h00;
            12'hFB1: q = 8'h00;
            12'hFB2: q = 8'h00;
            12'hFB3: q = 8'h00;
            12'hFB4: q = 8'h00;
            12'hFB5: q = 8'h00;
            12'hFB6: q = 8'h00;
            12'hFB7: q = 8'h00;
            12'hFB8: q = 8'h00;
            12'hFB9: q = 8'h00;
            12'hFBA: q = 8'h00;
            12'hFBB: q = 8'h00;
            12'hFBC: q = 8'h00;
            12'hFBD: q = 8'h00;
            12'hFBE: q = 8'h00;
            12'hFBF: q = 8'h00;
            12'hFC0: q = 8'h00;
            12'hFC1: q = 8'h00;
            12'hFC2: q = 8'h00;
            12'hFC3: q = 8'h00;
            12'hFC4: q = 8'h00;
            12'hFC5: q = 8'h00;
            12'hFC6: q = 8'h00;
            12'hFC7: q = 8'h00;
            12'hFC8: q = 8'h00;
            12'hFC9: q = 8'h00;
            12'hFCA: q = 8'h00;
            12'hFCB: q = 8'h00;
            12'hFCC: q = 8'h00;
            12'hFCD: q = 8'h00;
            12'hFCE: q = 8'h00;
            12'hFCF: q = 8'h00;
            12'hFD0: q = 8'h00;
            12'hFD1: q = 8'h00;
            12'hFD2: q = 8'h00;
            12'hFD3: q = 8'h00;
            12'hFD4: q = 8'h00;
            12'hFD5: q = 8'h00;
            12'hFD6: q = 8'h00;
            12'hFD7: q = 8'h00;
            12'hFD8: q = 8'h00;
            12'hFD9: q = 8'h00;
            12'hFDA: q = 8'h00;
            12'hFDB: q = 8'h00;
            12'hFDC: q = 8'h00;
            12'hFDD: q = 8'h00;
            12'hFDE: q = 8'h00;
            12'hFDF: q = 8'h00;
            12'hFE0: q = 8'h00;
            12'hFE1: q = 8'h00;
            12'hFE2: q = 8'h00;
            12'hFE3: q = 8'h00;
            12'hFE4: q = 8'h00;
            12'hFE5: q = 8'h00;
            12'hFE6: q = 8'h00;
            12'hFE7: q = 8'h00;
            12'hFE8: q = 8'h00;
            12'hFE9: q = 8'h00;
            12'hFEA: q = 8'h00;
            12'hFEB: q = 8'h00;
            12'hFEC: q = 8'h00;
            12'hFED: q = 8'h00;
            12'hFEE: q = 8'h00;
            12'hFEF: q = 8'h00;
            12'hFF0: q = 8'h00;
            12'hFF1: q = 8'h00;
            12'hFF2: q = 8'h00;
            12'hFF3: q = 8'h00;
            12'hFF4: q = 8'h00;
            12'hFF5: q = 8'h00;
            12'hFF6: q = 8'h00;
            12'hFF7: q = 8'h00;
            12'hFF8: q = 8'h00;
            12'hFF9: q = 8'h00;
            12'hFFA: q = 8'h00;
            12'hFFB: q = 8'h00;
            12'hFFC: q = 8'h00;
            12'hFFD: q = 8'h00;
            12'hFFE: q = 8'h00;
            12'hFFF: q = 8'h00;

			default:q = 0;
			
			
			
		endcase
		
endmodule
